 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT cap_mim 
+ C0_000 C1_000
+ C0_039 C1_039
+ C0_080 C1_080
+ C0_000 C1_000
+ C0_039 C1_039
+ C0_080 C1_080


C000 C0_000 C1_000 sky130_fd_pr__model__cap_mim AREA=4 PJ=8

C039 C0_039 C1_039 sky130_fd_pr__model__cap_mim AREA=1344 PJ=148

C080 C0_080 C1_080 sky130_fd_pr__model__cap_mim AREA=6724 PJ=328

C000 C0_000 C1_000 sky130_fd_pr__model__cap_mim_m4 AREA=4 PJ=8

C039 C0_039 C1_039 sky130_fd_pr__model__cap_mim_m4 AREA=1344 PJ=148

C080 C0_080 C1_080 sky130_fd_pr__model__cap_mim_m4 AREA=6724 PJ=328

.ENDS