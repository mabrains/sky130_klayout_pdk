 
* Copyright 2022 Mabrains
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Affero General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Affero General Public License for more details.
* 
* You should have received a copy of the GNU Affero General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.

.SUBCKT sky130_fd_pr__cap_vpp_02p7x41p1_m1m2m3m4_shieldl1_fingercap C0 C1 SUB

Cx C0 C1 SUB sky130_fd_pr__cap_vpp_02p7x41p1_m1m2m3m4_shieldl1_fingercap

.ENDS 
