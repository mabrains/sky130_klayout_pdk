 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT pfet BULK
+ SOURCE0 GATE0 DRAIN0
+ SOURCE31 GATE31 DRAIN31
+ SOURCE63 GATE63 DRAIN63
+ SOURCE0 GATE0 DRAIN0
+ SOURCE31 GATE31 DRAIN31
+ SOURCE63 GATE63 DRAIN63
+ SOURCE0 GATE0 DRAIN0
+ SOURCE31 GATE31 DRAIN31
+ SOURCE63 GATE63 DRAIN63
+ SOURCE0 GATE0 DRAIN0
+ SOURCE31 GATE31 DRAIN31
+ SOURCE63 GATE63 DRAIN63
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ DRAIN GATE SOURCE BULK
+ Bulk DRAIN GATE SOURCE
+ DRAIN GATE SOURCE BULK
+ 


M0 SOURCE0 GATE0 DRAIN0 BULK sky130_fd_pr__pfet_01v8 w=0.42 l=0.15 nf=1 

+ m=1 ad=0.9500400000000001 as=0.9500400000000001 pd=8.292000000000002 ps=8.292000000000002 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

+ m=1 ad=0.8526 as=0.8526 pd=9.94 ps=9.94 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

M0 SOURCE0 GATE0 DRAIN0 BULK sky130_fd_pr__pfet_01v8_hvt w=0.42 l=0.15 nf=1 

+ m=1 ad=0.9500400000000001 as=0.9500400000000001 pd=8.292000000000002 ps=8.292000000000002 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

+ m=1 ad=0.8526 as=0.8526 pd=9.94 ps=9.94 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

M0 SOURCE0 GATE0 DRAIN0 BULK sky130_fd_pr__pfet_01v8_lvt w=0.42 l=0.15 nf=1 

+ m=1 ad=0.9500400000000001 as=0.9500400000000001 pd=8.292000000000002 ps=8.292000000000002 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

+ m=1 ad=0.8526 as=0.8526 pd=9.94 ps=9.94 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

M0 SOURCE0 GATE0 DRAIN0 BULK sky130_fd_pr__pfet_g5v0d10v5 w=0.42 l=0.15 nf=1 

+ m=1 ad=0.9500400000000001 as=0.9500400000000001 pd=8.292000000000002 ps=8.292000000000002 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

+ m=1 ad=0.8526 as=0.8526 pd=9.94 ps=9.94 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF02W1p68L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF02W2p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF04W0p84L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF04W2p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF04W3p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF06W0p84L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF06W1p68L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF06W2p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF06W3p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF08W0p84L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aF08W1p68L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM02W1p65L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM02W1p65L0p18

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM02W1p65L0p25

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM02W3p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM02W3p00L0p18

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM02W3p00L0p25

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM02W5p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM02W5p00L0p18

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM02W5p00L0p25

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM04W1p65L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM04W1p65L0p18

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM04W1p65L0p25

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p18

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p25

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p18

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p25

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p18

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p25

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p18

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p25

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p18

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p25

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p18

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p25

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p18

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p25

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p18

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p25

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_hcM04W3p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_hcM04W5p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_lvt_aM02W3p00L0p35

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_lvt_aM02W3p00L0p50

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_lvt_aM02W5p00L0p35

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_lvt_aM02W5p00L0p50

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_lvt_aM04W3p00L0p35

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_lvt_aM04W3p00L0p50

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p35

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p50

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_mcM04W3p00L0p15

Mx Bulk DRAIN GATE SOURCE sky130_fd_pr__rf_pfet_01v8_mcM04W5p00L0p15

Mx DRAIN GATE SOURCE BULK sky130_fd_pr__rf_pfet_01v8_mvt_aF02W0p84L0p15

Mx  sky130_fd_pr__rf_pfet_20v0_withptap

.ENDS