* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hdll__mux2_16 A0 A1 S VGND VNB VPB VPWR X
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I X:O
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=4 w=0.65U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=4 w=0.65U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=4 w=0.65U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=4 w=0.65U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=2 w=0.65U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=16 w=0.65U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=4 w=1.0U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=4 w=1.0U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=4 w=1.0U l=0.18U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=4 w=1.0U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=2 w=1.0U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=16 w=1.0U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_hdll__mux2_16
