 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__model__cap_mim
+ C0_0 C1_0
+ C0_1 C1_1
+ C0_2 C1_2
+ C0_3 C1_3
+ C0_4 C1_4
+ C0_5 C1_5
+ C0_6 C1_6
+ C0_7 C1_7
+ C0_8 C1_8
+ C0_9 C1_9
+ C0_10 C1_10
+ C0_11 C1_11
+ C0_12 C1_12
+ C0_13 C1_13
+ C0_14 C1_14
+ C0_15 C1_15
+ C0_16 C1_16
+ C0_17 C1_17
+ C0_18 C1_18
+ C0_19 C1_19
+ C0_20 C1_20
+ C0_21 C1_21
+ C0_22 C1_22
+ C0_23 C1_23
+ C0_24 C1_24
+ C0_25 C1_25
+ C0_26 C1_26
+ C0_27 C1_27
+ C0_28 C1_28
+ C0_29 C1_29
+ C0_30 C1_30
+ C0_31 C1_31
+ C0_32 C1_32
+ C0_33 C1_33
+ C0_34 C1_34
+ C0_35 C1_35
+ C0_36 C1_36
+ C0_37 C1_37
+ C0_38 C1_38
+ C0_39 C1_39
+ C0_40 C1_40
+ C0_41 C1_41
+ C0_42 C1_42
+ C0_43 C1_43
+ C0_44 C1_44
+ C0_45 C1_45
+ C0_46 C1_46
+ C0_47 C1_47
+ C0_48 C1_48
+ C0_49 C1_49
+ C0_50 C1_50
+ C0_51 C1_51
+ C0_52 C1_52
+ C0_53 C1_53
+ C0_54 C1_54
+ C0_55 C1_55
+ C0_56 C1_56
+ C0_57 C1_57
+ C0_58 C1_58
+ C0_59 C1_59
+ C0_60 C1_60
+ C0_61 C1_61
+ C0_62 C1_62
+ C0_63 C1_63
+ C0_64 C1_64
+ C0_65 C1_65
+ C0_66 C1_66
+ C0_67 C1_67
+ C0_68 C1_68
+ C0_69 C1_69
+ C0_70 C1_70
+ C0_71 C1_71
+ C0_72 C1_72
+ C0_73 C1_73
+ C0_74 C1_74
+ C0_75 C1_75
+ C0_76 C1_76
+ C0_77 C1_77
+ C0_78 C1_78
+ C0_79 C1_79
+ C0_80 C1_80

C0 C0_0 C1_0 sky130_fd_pr__model__cap_mim AREA=4 PJ=8

C1 C0_1 C1_1 sky130_fd_pr__model__cap_mim AREA=24 PJ=28

C2 C0_2 C1_2 sky130_fd_pr__model__cap_mim AREA=44 PJ=48

C3 C0_3 C1_3 sky130_fd_pr__model__cap_mim AREA=64 PJ=68

C4 C0_4 C1_4 sky130_fd_pr__model__cap_mim AREA=84 PJ=88

C5 C0_5 C1_5 sky130_fd_pr__model__cap_mim AREA=104 PJ=108

C6 C0_6 C1_6 sky130_fd_pr__model__cap_mim AREA=124 PJ=128

C7 C0_7 C1_7 sky130_fd_pr__model__cap_mim AREA=144 PJ=148

C8 C0_8 C1_8 sky130_fd_pr__model__cap_mim AREA=164 PJ=168

C9 C0_9 C1_9 sky130_fd_pr__model__cap_mim AREA=24 PJ=28

C10 C0_10 C1_10 sky130_fd_pr__model__cap_mim AREA=144 PJ=48

C11 C0_11 C1_11 sky130_fd_pr__model__cap_mim AREA=264 PJ=68

C12 C0_12 C1_12 sky130_fd_pr__model__cap_mim AREA=384 PJ=88

C13 C0_13 C1_13 sky130_fd_pr__model__cap_mim AREA=504 PJ=108

C14 C0_14 C1_14 sky130_fd_pr__model__cap_mim AREA=624 PJ=128

C15 C0_15 C1_15 sky130_fd_pr__model__cap_mim AREA=744 PJ=148

C16 C0_16 C1_16 sky130_fd_pr__model__cap_mim AREA=864 PJ=168

C17 C0_17 C1_17 sky130_fd_pr__model__cap_mim AREA=984 PJ=188

C18 C0_18 C1_18 sky130_fd_pr__model__cap_mim AREA=44 PJ=48

C19 C0_19 C1_19 sky130_fd_pr__model__cap_mim AREA=264 PJ=68

C20 C0_20 C1_20 sky130_fd_pr__model__cap_mim AREA=484 PJ=88

C21 C0_21 C1_21 sky130_fd_pr__model__cap_mim AREA=704 PJ=108

C22 C0_22 C1_22 sky130_fd_pr__model__cap_mim AREA=924 PJ=128

C23 C0_23 C1_23 sky130_fd_pr__model__cap_mim AREA=1144 PJ=148

C24 C0_24 C1_24 sky130_fd_pr__model__cap_mim AREA=1364 PJ=168

C25 C0_25 C1_25 sky130_fd_pr__model__cap_mim AREA=1584 PJ=188

C26 C0_26 C1_26 sky130_fd_pr__model__cap_mim AREA=1804 PJ=208

C27 C0_27 C1_27 sky130_fd_pr__model__cap_mim AREA=64 PJ=68

C28 C0_28 C1_28 sky130_fd_pr__model__cap_mim AREA=384 PJ=88

C29 C0_29 C1_29 sky130_fd_pr__model__cap_mim AREA=704 PJ=108

C30 C0_30 C1_30 sky130_fd_pr__model__cap_mim AREA=1024 PJ=128

C31 C0_31 C1_31 sky130_fd_pr__model__cap_mim AREA=1344 PJ=148

C32 C0_32 C1_32 sky130_fd_pr__model__cap_mim AREA=1664 PJ=168

C33 C0_33 C1_33 sky130_fd_pr__model__cap_mim AREA=1984 PJ=188

C34 C0_34 C1_34 sky130_fd_pr__model__cap_mim AREA=2304 PJ=208

C35 C0_35 C1_35 sky130_fd_pr__model__cap_mim AREA=2624 PJ=228

C36 C0_36 C1_36 sky130_fd_pr__model__cap_mim AREA=84 PJ=88

C37 C0_37 C1_37 sky130_fd_pr__model__cap_mim AREA=504 PJ=108

C38 C0_38 C1_38 sky130_fd_pr__model__cap_mim AREA=924 PJ=128

C39 C0_39 C1_39 sky130_fd_pr__model__cap_mim AREA=1344 PJ=148

C40 C0_40 C1_40 sky130_fd_pr__model__cap_mim AREA=1764 PJ=168

C41 C0_41 C1_41 sky130_fd_pr__model__cap_mim AREA=2184 PJ=188

C42 C0_42 C1_42 sky130_fd_pr__model__cap_mim AREA=2604 PJ=208

C43 C0_43 C1_43 sky130_fd_pr__model__cap_mim AREA=3024 PJ=228

C44 C0_44 C1_44 sky130_fd_pr__model__cap_mim AREA=3444 PJ=248

C45 C0_45 C1_45 sky130_fd_pr__model__cap_mim AREA=104 PJ=108

C46 C0_46 C1_46 sky130_fd_pr__model__cap_mim AREA=624 PJ=128

C47 C0_47 C1_47 sky130_fd_pr__model__cap_mim AREA=1144 PJ=148

C48 C0_48 C1_48 sky130_fd_pr__model__cap_mim AREA=1664 PJ=168

C49 C0_49 C1_49 sky130_fd_pr__model__cap_mim AREA=2184 PJ=188

C50 C0_50 C1_50 sky130_fd_pr__model__cap_mim AREA=2704 PJ=208

C51 C0_51 C1_51 sky130_fd_pr__model__cap_mim AREA=3224 PJ=228

C52 C0_52 C1_52 sky130_fd_pr__model__cap_mim AREA=3744 PJ=248

C53 C0_53 C1_53 sky130_fd_pr__model__cap_mim AREA=4264 PJ=268

C54 C0_54 C1_54 sky130_fd_pr__model__cap_mim AREA=124 PJ=128

C55 C0_55 C1_55 sky130_fd_pr__model__cap_mim AREA=744 PJ=148

C56 C0_56 C1_56 sky130_fd_pr__model__cap_mim AREA=1364 PJ=168

C57 C0_57 C1_57 sky130_fd_pr__model__cap_mim AREA=1984 PJ=188

C58 C0_58 C1_58 sky130_fd_pr__model__cap_mim AREA=2604 PJ=208

C59 C0_59 C1_59 sky130_fd_pr__model__cap_mim AREA=3224 PJ=228

C60 C0_60 C1_60 sky130_fd_pr__model__cap_mim AREA=3844 PJ=248

C61 C0_61 C1_61 sky130_fd_pr__model__cap_mim AREA=4464 PJ=268

C62 C0_62 C1_62 sky130_fd_pr__model__cap_mim AREA=5084 PJ=288

C63 C0_63 C1_63 sky130_fd_pr__model__cap_mim AREA=144 PJ=148

C64 C0_64 C1_64 sky130_fd_pr__model__cap_mim AREA=864 PJ=168

C65 C0_65 C1_65 sky130_fd_pr__model__cap_mim AREA=1584 PJ=188

C66 C0_66 C1_66 sky130_fd_pr__model__cap_mim AREA=2304 PJ=208

C67 C0_67 C1_67 sky130_fd_pr__model__cap_mim AREA=3024 PJ=228

C68 C0_68 C1_68 sky130_fd_pr__model__cap_mim AREA=3744 PJ=248

C69 C0_69 C1_69 sky130_fd_pr__model__cap_mim AREA=4464 PJ=268

C70 C0_70 C1_70 sky130_fd_pr__model__cap_mim AREA=5184 PJ=288

C71 C0_71 C1_71 sky130_fd_pr__model__cap_mim AREA=5904 PJ=308

C72 C0_72 C1_72 sky130_fd_pr__model__cap_mim AREA=164 PJ=168

C73 C0_73 C1_73 sky130_fd_pr__model__cap_mim AREA=984 PJ=188

C74 C0_74 C1_74 sky130_fd_pr__model__cap_mim AREA=1804 PJ=208

C75 C0_75 C1_75 sky130_fd_pr__model__cap_mim AREA=2624 PJ=228

C76 C0_76 C1_76 sky130_fd_pr__model__cap_mim AREA=3444 PJ=248

C77 C0_77 C1_77 sky130_fd_pr__model__cap_mim AREA=4264 PJ=268

C78 C0_78 C1_78 sky130_fd_pr__model__cap_mim AREA=5084 PJ=288

C79 C0_79 C1_79 sky130_fd_pr__model__cap_mim AREA=5904 PJ=308

C80 C0_80 C1_80 sky130_fd_pr__model__cap_mim AREA=6724 PJ=328

.ENDS