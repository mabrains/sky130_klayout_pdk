*** HVL Include files.

.include ./hvl_cdl/sky130_fd_sc_hvl__a21o_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__a21oi_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__a22o_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__a22oi_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__and2_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__and3_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__buf_16.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__buf_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__buf_2.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__buf_32.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__buf_4.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__buf_8.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__decap_4.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__decap_8.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__dfrbp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__dfrtp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__dfsbp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__dfstp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__dfxbp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__dfxtp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__dlclkp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__dlrtp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__dlxtp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__einvn_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__einvp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__inv_16.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__inv_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__inv_2.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__inv_4.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__inv_8.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__lsbufhv2hv_hl_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__lsbufhv2hv_lh_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__lsbufhv2lv_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__lsbufhv2lv_simple_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__lsbuflv2hv_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__mux2_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__mux4_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__nand2_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__nand3_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__nor2_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__nor3_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__o21a_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__o21ai_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__o22a_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__o22ai_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__or2_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__or3_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__probec_p_8.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__probe_p_8.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__schmittbuf_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__sdfrbp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__sdfrtp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__sdfsbp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__sdfstp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__sdfxbp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__sdfxtp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__sdlclkp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__sdlxtp_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__xnor2_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__xor2_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__conb_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__diode_2.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__fill_1.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__fill_2.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__fill_4.cdl
.include ./hvl_cdl/sky130_fd_sc_hvl__fill_8.cdl
