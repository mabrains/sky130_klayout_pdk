 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__diode_pw2nd_05v5_lvt
+ D0_0 D1_0
+ D0_1 D1_1
+ D0_2 D1_2
+ D0_3 D1_3
+ D0_4 D1_4
+ D0_5 D1_5
+ D0_6 D1_6
+ D0_7 D1_7
+ D0_8 D1_8
+ D0_9 D1_9
+ D0_10 D1_10
+ D0_11 D1_11
+ D0_12 D1_12
+ D0_13 D1_13
+ D0_14 D1_14
+ D0_15 D1_15
+ D0_16 D1_16
+ D0_17 D1_17
+ D0_18 D1_18
+ D0_19 D1_19
+ D0_20 D1_20
+ D0_21 D1_21
+ D0_22 D1_22
+ D0_23 D1_23
+ D0_24 D1_24
+ D0_25 D1_25
+ D0_26 D1_26
+ D0_27 D1_27
+ D0_28 D1_28
+ D0_29 D1_29
+ D0_30 D1_30
+ D0_31 D1_31
+ D0_32 D1_32
+ D0_33 D1_33
+ D0_34 D1_34
+ D0_35 D1_35
+ D0_36 D1_36
+ D0_37 D1_37
+ D0_38 D1_38
+ D0_39 D1_39
+ D0_40 D1_40
+ D0_41 D1_41
+ D0_42 D1_42
+ D0_43 D1_43
+ D0_44 D1_44
+ D0_45 D1_45
+ D0_46 D1_46
+ D0_47 D1_47
+ D0_48 D1_48
+ D0_49 D1_49
+ D0_50 D1_50
+ D0_51 D1_51
+ D0_52 D1_52
+ D0_53 D1_53
+ D0_54 D1_54
+ D0_55 D1_55
+ D0_56 D1_56
+ D0_57 D1_57
+ D0_58 D1_58
+ D0_59 D1_59
+ D0_60 D1_60
+ D0_61 D1_61
+ D0_62 D1_62
+ D0_63 D1_63

D0 D0_0 D1_0 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=0.2 PJ=1.8

D1 D0_1 D1_1 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=0.41 PJ=2.7

D2 D0_2 D1_2 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=0.61 PJ=3.6

D3 D0_3 D1_3 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=0.81 PJ=4.5

D4 D0_4 D1_4 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=1.01 PJ=5.4

D5 D0_5 D1_5 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=1.22 PJ=6.3

D6 D0_6 D1_6 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=1.42 PJ=7.2

D7 D0_7 D1_7 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=1.62 PJ=8.1

D8 D0_8 D1_8 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=0.41 PJ=2.7

D9 D0_9 D1_9 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=0.81 PJ=3.6

D10 D0_10 D1_10 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=1.22 PJ=4.5

D11 D0_11 D1_11 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=1.62 PJ=5.4

D12 D0_12 D1_12 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=2.02 PJ=6.3

D13 D0_13 D1_13 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=2.43 PJ=7.2

D14 D0_14 D1_14 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=2.84 PJ=8.1

D15 D0_15 D1_15 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=3.24 PJ=9.0

D16 D0_16 D1_16 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=0.61 PJ=3.6

D17 D0_17 D1_17 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=1.22 PJ=4.5

D18 D0_18 D1_18 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=1.82 PJ=5.4

D19 D0_19 D1_19 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=2.43 PJ=6.3

D20 D0_20 D1_20 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=3.04 PJ=7.2

D21 D0_21 D1_21 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=3.65 PJ=8.1

D22 D0_22 D1_22 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=4.25 PJ=9.0

D23 D0_23 D1_23 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=4.86 PJ=9.9

D24 D0_24 D1_24 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=0.81 PJ=4.5

D25 D0_25 D1_25 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=1.62 PJ=5.4

D26 D0_26 D1_26 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=2.43 PJ=6.3

D27 D0_27 D1_27 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=3.24 PJ=7.2

D28 D0_28 D1_28 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=4.05 PJ=8.1

D29 D0_29 D1_29 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=4.86 PJ=9.0

D30 D0_30 D1_30 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=5.67 PJ=9.9

D31 D0_31 D1_31 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=6.48 PJ=10.8

D32 D0_32 D1_32 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=1.01 PJ=5.4

D33 D0_33 D1_33 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=2.02 PJ=6.3

D34 D0_34 D1_34 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=3.04 PJ=7.2

D35 D0_35 D1_35 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=4.05 PJ=8.1

D36 D0_36 D1_36 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=5.06 PJ=9.0

D37 D0_37 D1_37 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=6.08 PJ=9.9

D38 D0_38 D1_38 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=7.09 PJ=10.8

D39 D0_39 D1_39 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=8.1 PJ=11.7

D40 D0_40 D1_40 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=1.22 PJ=6.3

D41 D0_41 D1_41 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=2.43 PJ=7.2

D42 D0_42 D1_42 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=3.65 PJ=8.1

D43 D0_43 D1_43 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=4.86 PJ=9.0

D44 D0_44 D1_44 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=6.08 PJ=9.9

D45 D0_45 D1_45 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=7.29 PJ=10.8

D46 D0_46 D1_46 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=8.51 PJ=11.7

D47 D0_47 D1_47 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=9.72 PJ=12.6

D48 D0_48 D1_48 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=1.42 PJ=7.2

D49 D0_49 D1_49 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=2.84 PJ=8.1

D50 D0_50 D1_50 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=4.25 PJ=9.0

D51 D0_51 D1_51 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=5.67 PJ=9.9

D52 D0_52 D1_52 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=7.09 PJ=10.8

D53 D0_53 D1_53 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=8.51 PJ=11.7

D54 D0_54 D1_54 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=9.92 PJ=12.6

D55 D0_55 D1_55 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=11.34 PJ=13.5

D56 D0_56 D1_56 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=1.62 PJ=8.1

D57 D0_57 D1_57 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=3.24 PJ=9.0

D58 D0_58 D1_58 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=4.86 PJ=9.9

D59 D0_59 D1_59 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=6.48 PJ=10.8

D60 D0_60 D1_60 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=8.1 PJ=11.7

D61 D0_61 D1_61 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=9.72 PJ=12.6

D62 D0_62 D1_62 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=11.34 PJ=13.5

D63 D0_63 D1_63 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=12.96 PJ=14.4

.ENDS