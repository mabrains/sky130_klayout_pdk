 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT nfet SUBSTRATE
+ SOURCE0 GATE0 DRAIN0
+ SOURCE31 GATE31 DRAIN31
+ SOURCE63 GATE63 DRAIN63
+ SOURCE0 GATE0 DRAIN0
+ SOURCE31 GATE31 DRAIN31
+ SOURCE63 GATE63 DRAIN63
+ SOURCE0 GATE0 DRAIN0
+ SOURCE31 GATE31 DRAIN31
+ SOURCE63 GATE63 DRAIN63
+ SOURCE0 GATE0 DRAIN0
+ SOURCE31 GATE31 DRAIN31
+ SOURCE63 GATE63 DRAIN63
+ SOURCE0 GATE0 DRAIN0
+ SOURCE31 GATE31 DRAIN31
+ SOURCE63 GATE63 DRAIN63
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ GATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ 
+ 
+ D PSUB S
+ 
+ D G PSUB S
+ 
+ 
+ 
+ D PSUB S
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE
+ DRAIN GATE SOURCE SUBSTRATE


M0 SOURCE0 GATE0 DRAIN0 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=0.15 nf=1 

+ m=1 ad=0.9500400000000001 as=0.9500400000000001 pd=8.292000000000002 ps=8.292000000000002 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

+ m=1 ad=0.8526 as=0.8526 pd=9.94 ps=9.94 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

M0 SOURCE0 GATE0 DRAIN0 SUBSTRATE sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15 nf=1 

+ m=1 ad=0.9500400000000001 as=0.9500400000000001 pd=8.292000000000002 ps=8.292000000000002 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

+ m=1 ad=0.8526 as=0.8526 pd=9.94 ps=9.94 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

M0 SOURCE0 GATE0 DRAIN0 SUBSTRATE sky130_fd_pr__nfet_03v3_nvt w=0.42 l=0.15 nf=1 

+ m=1 ad=0.9500400000000001 as=0.9500400000000001 pd=8.292000000000002 ps=8.292000000000002 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

+ m=1 ad=0.8526 as=0.8526 pd=9.94 ps=9.94 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

M0 SOURCE0 GATE0 DRAIN0 SUBSTRATE sky130_fd_pr__nfet_05v0_nvt w=0.42 l=0.15 nf=1 

+ m=1 ad=0.9500400000000001 as=0.9500400000000001 pd=8.292000000000002 ps=8.292000000000002 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

+ m=1 ad=0.8526 as=0.8526 pd=9.94 ps=9.94 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

M0 SOURCE0 GATE0 DRAIN0 SUBSTRATE sky130_fd_pr__nfet_g5v0d10v5 w=0.42 l=0.15 nf=1 

+ m=1 ad=0.9500400000000001 as=0.9500400000000001 pd=8.292000000000002 ps=8.292000000000002 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

+ m=1 ad=0.8526 as=0.8526 pd=9.94 ps=9.94 nrd=0.0531135531135531 nrs=0.0531135531135531 sa=0 sb=0 sd=0

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W3p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W3p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM04W1p65L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM04W1p65L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM04W1p65L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM04W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM04W3p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM04W3p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_hcM04W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_hcM04W5p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p84L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF02W1p65L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF02W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p42L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF04W1p65L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF04W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF06W0p42L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF06W0p84L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF06W1p65L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF06W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF08W0p42L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF08W0p84L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF08W1p65L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM02W1p65L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM02W1p65L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM02W1p65L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM02W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM02W3p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM02W3p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p18

Mx GATE sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM04W1p65L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM04W1p65L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM04W1p65L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM04W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM04W3p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM04W3p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM02W1p65L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM02W1p65L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM02W1p65L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM02W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM02W3p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM02W3p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM02W5p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM02W5p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM02W5p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM04W1p65L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM04W1p65L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM04W1p65L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM04W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM04W3p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM04W3p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM04W5p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM04W5p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM04W5p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM02W1p65L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM02W1p65L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM02W1p65L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM02W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM02W3p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM02W3p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM02W5p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM02W5p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM02W5p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM04W1p65L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM04W1p65L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM04W1p65L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM04W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM04W3p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM04W3p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM04W5p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM04W5p00L0p18

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_cM04W5p00L0p25

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_mcM04W3p00L0p15

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_mcM04W5p00L0p15

Mx  sky130_fd_pr__rf_nfet_20v0_aup

Mx  sky130_fd_pr__rf_nfet_20v0_noptap_iso

Mx D PSUB S sky130_fd_pr__rf_nfet_20v0_nvt_aup

Mx  sky130_fd_pr__rf_nfet_20v0_nvt_noptap_iso

Mx D G PSUB S sky130_fd_pr__rf_nfet_20v0_nvt_withptap

Mx  sky130_fd_pr__rf_nfet_20v0_nvt_withptap_iso

Mx  sky130_fd_pr__rf_nfet_20v0_withptap

Mx  sky130_fd_pr__rf_nfet_20v0_withptap_iso

Mx D PSUB S sky130_fd_pr__rf_nfet_20v0_zvt_withptap

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W3p00L0p50

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W5p00L0p50

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W7p00L0p50

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W3p00L0p50

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W5p00L0p50

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W7p00L0p50

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W3p00L0p50

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W5p00L0p50

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W3p00L0p50

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00L0p50

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00L0p50

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W3p00L0p50

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W5p00L0p50

Mx DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00L0p50

.ENDS