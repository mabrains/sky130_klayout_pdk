 
* Copyright 2022 Mabrains
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Affero General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Affero General Public License for more details.
* 
* You should have received a copy of the GNU Affero General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM04W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE

Mx_dim_fail DRAIN_dim_fail GATE_dim_fail SOURCE_dim_fail SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM04W1p65L0p18 w=6.6u l=0.18u nf=4 m=1 ad=0.2392p as=0.2392p pd=2.81u ps=2.81u nrd=0.1758 nrs=0.1758 sa=0 sb=0 sd=0

.ENDS