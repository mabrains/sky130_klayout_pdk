 
* Copyright 2022 Mabrains
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Affero General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Affero General Public License for more details.
* 
* You should have received a copy of the GNU Affero General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.

.SUBCKT sky130_fd_pr__cap_var_lvt SUBSTRATE
+ C0_000 C1_000
+ C0_001 C1_001
+ C0_002 C1_002
+ C0_003 C1_003
+ C0_004 C1_004
+ C0_005 C1_005
+ C0_006 C1_006
+ C0_007 C1_007
+ C0_008 C1_008
+ C0_009 C1_009
+ C0_010 C1_010
+ C0_011 C1_011
+ C0_012 C1_012
+ C0_013 C1_013
+ C0_014 C1_014
+ C0_015 C1_015
+ C0_016 C1_016
+ C0_017 C1_017
+ C0_018 C1_018
+ C0_019 C1_019
+ C0_020 C1_020
+ C0_021 C1_021
+ C0_022 C1_022
+ C0_023 C1_023
+ C0_024 C1_024
+ C0_025 C1_025
+ C0_026 C1_026
+ C0_027 C1_027
+ C0_028 C1_028
+ C0_029 C1_029
+ C0_030 C1_030
+ C0_031 C1_031
+ C0_032 C1_032
+ C0_033 C1_033
+ C0_034 C1_034
+ C0_035 C1_035
+ C0_036 C1_036
+ C0_037 C1_037
+ C0_038 C1_038
+ C0_039 C1_039
+ C0_040 C1_040
+ C0_041 C1_041
+ C0_042 C1_042
+ C0_043 C1_043
+ C0_044 C1_044
+ C0_045 C1_045
+ C0_046 C1_046
+ C0_047 C1_047
+ C0_048 C1_048
+ C0_049 C1_049
+ C0_050 C1_050
+ C0_051 C1_051
+ C0_052 C1_052
+ C0_053 C1_053
+ C0_054 C1_054
+ C0_055 C1_055
+ C0_056 C1_056
+ C0_057 C1_057
+ C0_058 C1_058
+ C0_059 C1_059
+ C0_060 C1_060
+ C0_061 C1_061
+ C0_062 C1_062
+ C0_063 C1_063

C000 C0_000 C1_000 SUBSTRATE sky130_fd_pr__cap_var_lvt A=0.18p P=2.36u

C001 C0_001 C1_001 SUBSTRATE sky130_fd_pr__cap_var_lvt A=0.36p P=4.36u

C002 C0_002 C1_002 SUBSTRATE sky130_fd_pr__cap_var_lvt A=0.54p P=6.36u

C003 C0_003 C1_003 SUBSTRATE sky130_fd_pr__cap_var_lvt A=0.72p P=8.36u

C004 C0_004 C1_004 SUBSTRATE sky130_fd_pr__cap_var_lvt A=0.36p P=2.72u

C005 C0_005 C1_005 SUBSTRATE sky130_fd_pr__cap_var_lvt A=0.72p P=4.72u

C006 C0_006 C1_006 SUBSTRATE sky130_fd_pr__cap_var_lvt A=1.08p P=6.72u

C007 C0_007 C1_007 SUBSTRATE sky130_fd_pr__cap_var_lvt A=1.44p P=8.72u

C008 C0_008 C1_008 SUBSTRATE sky130_fd_pr__cap_var_lvt A=0.54p P=3.08u

C009 C0_009 C1_009 SUBSTRATE sky130_fd_pr__cap_var_lvt A=1.08p P=5.08u

C010 C0_010 C1_010 SUBSTRATE sky130_fd_pr__cap_var_lvt A=1.62p P=7.08u

C011 C0_011 C1_011 SUBSTRATE sky130_fd_pr__cap_var_lvt A=2.16p P=9.08u

C012 C0_012 C1_012 SUBSTRATE sky130_fd_pr__cap_var_lvt A=0.72p P=3.44u

C013 C0_013 C1_013 SUBSTRATE sky130_fd_pr__cap_var_lvt A=1.44p P=5.44u

C014 C0_014 C1_014 SUBSTRATE sky130_fd_pr__cap_var_lvt A=2.16p P=7.44u

C015 C0_015 C1_015 SUBSTRATE sky130_fd_pr__cap_var_lvt A=2.88p P=9.44u

C016 C0_016 C1_016 SUBSTRATE sky130_fd_pr__cap_var_lvt A=0.9p P=11.8u

C017 C0_017 C1_017 SUBSTRATE sky130_fd_pr__cap_var_lvt A=1.8p P=21.8u

C018 C0_018 C1_018 SUBSTRATE sky130_fd_pr__cap_var_lvt A=2.7p P=31.8u

C019 C0_019 C1_019 SUBSTRATE sky130_fd_pr__cap_var_lvt A=3.6p P=41.8u

C020 C0_020 C1_020 SUBSTRATE sky130_fd_pr__cap_var_lvt A=1.8p P=13.6u

C021 C0_021 C1_021 SUBSTRATE sky130_fd_pr__cap_var_lvt A=3.6p P=23.6u

C022 C0_022 C1_022 SUBSTRATE sky130_fd_pr__cap_var_lvt A=5.4p P=33.6u

C023 C0_023 C1_023 SUBSTRATE sky130_fd_pr__cap_var_lvt A=7.2p P=43.6u

C024 C0_024 C1_024 SUBSTRATE sky130_fd_pr__cap_var_lvt A=2.7p P=15.4u

C025 C0_025 C1_025 SUBSTRATE sky130_fd_pr__cap_var_lvt A=5.4p P=25.4u

C026 C0_026 C1_026 SUBSTRATE sky130_fd_pr__cap_var_lvt A=8.1p P=35.4u

C027 C0_027 C1_027 SUBSTRATE sky130_fd_pr__cap_var_lvt A=10.8p P=45.4u

C028 C0_028 C1_028 SUBSTRATE sky130_fd_pr__cap_var_lvt A=3.6p P=17.2u

C029 C0_029 C1_029 SUBSTRATE sky130_fd_pr__cap_var_lvt A=7.2p P=27.2u

C030 C0_030 C1_030 SUBSTRATE sky130_fd_pr__cap_var_lvt A=10.8p P=37.2u

C031 C0_031 C1_031 SUBSTRATE sky130_fd_pr__cap_var_lvt A=14.4p P=47.2u

C032 C0_032 C1_032 SUBSTRATE sky130_fd_pr__cap_var_lvt A=1.62p P=21.24u

C033 C0_033 C1_033 SUBSTRATE sky130_fd_pr__cap_var_lvt A=3.24p P=39.24u

C034 C0_034 C1_034 SUBSTRATE sky130_fd_pr__cap_var_lvt A=4.86p P=57.24u

C035 C0_035 C1_035 SUBSTRATE sky130_fd_pr__cap_var_lvt A=6.48p P=75.24u

C036 C0_036 C1_036 SUBSTRATE sky130_fd_pr__cap_var_lvt A=3.24p P=24.48u

C037 C0_037 C1_037 SUBSTRATE sky130_fd_pr__cap_var_lvt A=6.48p P=42.48u

C038 C0_038 C1_038 SUBSTRATE sky130_fd_pr__cap_var_lvt A=9.72p P=60.48u

C039 C0_039 C1_039 SUBSTRATE sky130_fd_pr__cap_var_lvt A=12.96p P=78.48u

C040 C0_040 C1_040 SUBSTRATE sky130_fd_pr__cap_var_lvt A=4.86p P=27.72u

C041 C0_041 C1_041 SUBSTRATE sky130_fd_pr__cap_var_lvt A=9.72p P=45.72u

C042 C0_042 C1_042 SUBSTRATE sky130_fd_pr__cap_var_lvt A=14.58p P=63.72u

C043 C0_043 C1_043 SUBSTRATE sky130_fd_pr__cap_var_lvt A=19.44p P=81.72u

C044 C0_044 C1_044 SUBSTRATE sky130_fd_pr__cap_var_lvt A=6.48p P=30.96u

C045 C0_045 C1_045 SUBSTRATE sky130_fd_pr__cap_var_lvt A=12.96p P=48.96u

C046 C0_046 C1_046 SUBSTRATE sky130_fd_pr__cap_var_lvt A=19.44p P=66.96u

C047 C0_047 C1_047 SUBSTRATE sky130_fd_pr__cap_var_lvt A=25.92p P=84.96u

C048 C0_048 C1_048 SUBSTRATE sky130_fd_pr__cap_var_lvt A=2.34p P=30.68u

C049 C0_049 C1_049 SUBSTRATE sky130_fd_pr__cap_var_lvt A=4.68p P=56.68u

C050 C0_050 C1_050 SUBSTRATE sky130_fd_pr__cap_var_lvt A=7.02p P=82.68u

C051 C0_051 C1_051 SUBSTRATE sky130_fd_pr__cap_var_lvt A=9.36p P=108.68u

C052 C0_052 C1_052 SUBSTRATE sky130_fd_pr__cap_var_lvt A=4.68p P=35.36u

C053 C0_053 C1_053 SUBSTRATE sky130_fd_pr__cap_var_lvt A=9.36p P=61.36u

C054 C0_054 C1_054 SUBSTRATE sky130_fd_pr__cap_var_lvt A=14.04p P=87.36u

C055 C0_055 C1_055 SUBSTRATE sky130_fd_pr__cap_var_lvt A=18.72p P=113.36u

C056 C0_056 C1_056 SUBSTRATE sky130_fd_pr__cap_var_lvt A=7.02p P=40.04u

C057 C0_057 C1_057 SUBSTRATE sky130_fd_pr__cap_var_lvt A=14.04p P=66.04u

C058 C0_058 C1_058 SUBSTRATE sky130_fd_pr__cap_var_lvt A=21.06p P=92.04u

C059 C0_059 C1_059 SUBSTRATE sky130_fd_pr__cap_var_lvt A=28.08p P=118.04u

C060 C0_060 C1_060 SUBSTRATE sky130_fd_pr__cap_var_lvt A=9.36p P=44.72u

C061 C0_061 C1_061 SUBSTRATE sky130_fd_pr__cap_var_lvt A=18.72p P=70.72u

C062 C0_062 C1_062 SUBSTRATE sky130_fd_pr__cap_var_lvt A=28.08p P=96.72u

C063 C0_063 C1_063 SUBSTRATE sky130_fd_pr__cap_var_lvt A=37.44p P=122.72u

.ENDS