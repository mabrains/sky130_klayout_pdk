 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_20v0_nvt_aup D PSUB S

Mx D PSUB S sky130_fd_pr__rf_nfet_20v0_nvt_aup

Mx_net_fail D_net_fail PSUB S_net_fail sky130_fd_pr__rf_nfet_20v0_nvt_aup

Mx_dim_fail D_dim_fail PSUB S_dim_fail sky130_fd_pr__rf_nfet_20v0_nvt_aup

.ENDS