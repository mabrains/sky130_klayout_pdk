*** HDLL Include files.

.include ./hdll_cdl/sky130_fd_sc_hdll__a211o_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a211o_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a211oi_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a211oi_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a21bo_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a21bo_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a21boi_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a21boi_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a21o_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a21o_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a21oi_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a21oi_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a221oi_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a221oi_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a221oi_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a222oi_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a22o_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a22o_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a22o_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a22oi_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a22oi_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a22oi_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a2bb2o_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a2bb2o_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a2bb2o_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a2bb2oi_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a2bb2oi_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a2bb2oi_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a31o_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a31o_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a31oi_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a31oi_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a31oi_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a32o_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a32o_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a32o_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a32oi_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a32oi_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a32oi_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and2_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and2_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and2_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and2b_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and2b_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and2b_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and3_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and3_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and3_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and3b_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and3b_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and3b_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and4_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and4_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and4_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and4b_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and4b_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and4b_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and4bb_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and4bb_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and4bb_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__buf_12.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__buf_16.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__buf_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__buf_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__buf_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__buf_6.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__buf_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__bufbuf_16.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__bufbuf_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__bufinv_16.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__bufinv_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkbuf_12.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkbuf_16.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkbuf_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkbuf_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkbuf_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkbuf_6.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkbuf_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkinv_12.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkinv_16.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkinv_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkinv_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkinv_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkinv_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkinvlp_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkinvlp_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkmux2_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkmux2_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__clkmux2_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__decap_12.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__decap_3.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__decap_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__decap_6.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__decap_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dfrtp_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dfrtp_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dfrtp_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dfstp_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dfstp_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dfstp_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dlrtn_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dlrtn_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dlrtn_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dlrtp_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dlrtp_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dlrtp_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dlxtn_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dlxtn_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dlxtn_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dlygate4sd1_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dlygate4sd2_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__dlygate4sd3_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__ebufn_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__ebufn_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__ebufn_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__ebufn_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__einvn_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__einvn_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__einvn_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__einvn_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__einvp_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__einvp_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__einvp_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__einvp_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__inputiso0n_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__inputiso0p_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__inputiso1n_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__inputiso1p_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__inv_12.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__inv_16.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__inv_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__inv_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__inv_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__inv_6.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__inv_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__isobufsrc_16.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__isobufsrc_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__isobufsrc_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__isobufsrc_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__isobufsrc_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__mux2_12.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__mux2_16.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__mux2_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__mux2_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__mux2_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__mux2_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__mux2i_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__mux2i_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__mux2i_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__muxb16to1_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__muxb16to1_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__muxb16to1_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__muxb4to1_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__muxb4to1_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__muxb4to1_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__muxb8to1_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__muxb8to1_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__muxb8to1_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand2_12.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand2_16.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand2_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand2_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand2_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand2_6.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand2_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand2b_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand2b_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand2b_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand3_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand3_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand3_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand3b_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand3b_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand3b_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand4_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand4_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand4_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand4b_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand4b_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand4b_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand4bb_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand4bb_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nand4bb_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor2_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor2_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor2_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor2_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor2b_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor2b_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor2b_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor3_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor3_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor3_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor3b_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor3b_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor3b_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor4_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor4_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor4_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor4_6.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor4_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor4b_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor4b_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor4b_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor4bb_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor4bb_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__nor4bb_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o211a_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o211a_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o211ai_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o211ai_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o21a_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o21a_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o21ai_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o21ai_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o21ai_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o21ba_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o21ba_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o21ba_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o21bai_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o21bai_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o21bai_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o221a_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o221a_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o221a_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o221ai_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o221ai_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o221ai_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o22a_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o22a_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o22a_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o22ai_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o22ai_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o22ai_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o2bb2a_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o2bb2a_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o2bb2a_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o2bb2ai_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o2bb2ai_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o2bb2ai_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o31ai_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o31ai_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o31ai_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o32ai_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o32ai_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o32ai_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or2_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or2_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or2_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or2_6.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or2_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or2b_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or2b_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or2b_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or3_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or3_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or3_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or3b_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or3b_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or3b_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or4_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or4_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or4_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or4b_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or4b_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or4b_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or4bb_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or4bb_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__or4bb_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__probec_p_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__probe_p_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfbbp_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfrbp_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfrbp_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfrtn_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfrtp_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfrtp_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfrtp_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfsbp_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfsbp_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfstp_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfstp_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfstp_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfxbp_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfxbp_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfxtp_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfxtp_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdfxtp_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdlclkp_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdlclkp_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sdlclkp_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sedfxbp_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__sedfxbp_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__xnor2_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__xnor2_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__xnor2_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__xnor3_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__xnor3_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__xnor3_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__xor2_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__xor2_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__xor2_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__xor3_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__xor3_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__xor3_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a211o_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a211oi_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a21bo_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a21boi_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a21o_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a21o_6.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a21o_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a21oi_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__a31o_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and2_6.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__and2_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__conb_1.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__diode_2.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__diode_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__diode_6.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__diode_8.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o211a_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o211ai_4.cdl
.include ./hdll_cdl/sky130_fd_sc_hdll__o21a_4.cdl
