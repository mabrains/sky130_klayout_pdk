* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN2 X y VGND VNB nfet_01v8_lvt m=4 w=0.74U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8_lvt m=1 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8_lvt m=1 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8_lvt m=2 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8_lvt m=2 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8_lvt m=2 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8 m=4 w=1.12U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8 m=1 w=0.84U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8 m=1 w=0.84U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8 m=2 w=1.0U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8 m=2 w=1.0U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8 m=2 w=0.84U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_hs__o2bb2a_4
