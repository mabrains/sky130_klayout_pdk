* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hdll__nor2_8 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMP1 sndPA B Y VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65U l=0.15U mult=1 sa=0.265 sb=0.265
+ sd=0.28 area=0.063 perim=1.14
MMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65U l=0.15U mult=1 sa=0.265 sb=0.265
+ sd=0.28 area=0.063 perim=1.14
.ENDS sky130_fd_sc_hdll__nor2_8
