* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__schmittbuf_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
rI39 net069 VGND VNB sky130_fd_pr__res_generic_nd_hv m=1 w=0.29U l=1.355U
rI38 VPWR net32 VPB sky130_fd_pr__res_generic_pd_hv m=1 w=0.29U l=3.11U
MI5 net32 net36 net40 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MMN0 net36 A net40 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMN1 net40 A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMIN1 X net36 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI6 net069 net36 net56 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MMP0 VPWR A net56 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMP1 net56 A net36 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMIP1 X net36 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
.ENDS sky130_fd_sc_hvl__schmittbuf_1
