* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_lp__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net175 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net175 VPWR VPB pfet_01v8_hvt m=2 w=1.26U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N S0 VPWR VPB pfet_01v8_hvt m=2 w=1.26U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net110 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net110 VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net102 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net102 VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net90 VPB pfet_01v8_hvt m=1 w=0.84U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net90 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net203 VNB nfet_01v8 m=1 w=0.64U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net223 S1 net167 VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net214 VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net210 VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net214 M1 VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net203 M0 VGND VNB nfet_01v8 m=1 w=0.64U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net223 VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N S0 VGND VNB nfet_01v8 m=2 w=0.84U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net210 SET_B VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net175 S0 VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net167 SET_B VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net175 VGND VNB nfet_01v8 m=2 w=0.84U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS sky130_fd_sc_lp__sdfsbp_2
