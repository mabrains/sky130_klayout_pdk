* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or2b_1 A B_N VGND VNB VPB VPWR X
*.PININFO A:I B_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8 m=1 w=1.0U l=0.15U mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8 m=1 w=0.84U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8 m=1 w=1.12U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.55U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.55U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8_lvt m=1 w=0.55U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8_lvt m=1 w=0.74U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_hs__or2b_1
