* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_lp__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.26U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.26U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.26U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.26U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.84U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.84U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.84U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.84U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_lp__o211ai_4
