 
* Copyright 2022 Mabrains
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Affero General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Affero General Public License for more details.
* 
* You should have received a copy of the GNU Affero General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.

.SUBCKT sky130_fd_pr__cap_var_hvt SUBSTRATE
+ C0_000_net_fail C1_000_net_fail
+ C0_001_net_fail C1_001_net_fail
+ C0_002_net_fail C1_002_net_fail
+ C0_003_net_fail C1_003_net_fail
+ C0_004_net_fail C1_004_net_fail
+ C0_005_net_fail C1_005_net_fail
+ C0_006_net_fail C1_006_net_fail
+ C0_007_net_fail C1_007_net_fail
+ C0_008_net_fail C1_008_net_fail
+ C0_009_net_fail C1_009_net_fail
+ C0_010_net_fail C1_010_net_fail
+ C0_011_net_fail C1_011_net_fail
+ C0_012_net_fail C1_012_net_fail
+ C0_013_net_fail C1_013_net_fail
+ C0_014_net_fail C1_014_net_fail
+ C0_015_net_fail C1_015_net_fail
+ C0_016_net_fail C1_016_net_fail
+ C0_017_net_fail C1_017_net_fail
+ C0_018_net_fail C1_018_net_fail
+ C0_019_net_fail C1_019_net_fail
+ C0_020_net_fail C1_020_net_fail
+ C0_021_net_fail C1_021_net_fail
+ C0_022_net_fail C1_022_net_fail
+ C0_023_net_fail C1_023_net_fail
+ C0_024_net_fail C1_024_net_fail
+ C0_025_net_fail C1_025_net_fail
+ C0_026_net_fail C1_026_net_fail
+ C0_027_net_fail C1_027_net_fail
+ C0_028_net_fail C1_028_net_fail
+ C0_029_net_fail C1_029_net_fail
+ C0_030_net_fail C1_030_net_fail
+ C0_031_net_fail C1_031_net_fail
+ C0_032_net_fail C1_032_net_fail
+ C0_033_net_fail C1_033_net_fail
+ C0_034_net_fail C1_034_net_fail
+ C0_035_net_fail C1_035_net_fail
+ C0_036_net_fail C1_036_net_fail
+ C0_037_net_fail C1_037_net_fail
+ C0_038_net_fail C1_038_net_fail
+ C0_039_net_fail C1_039_net_fail
+ C0_040_net_fail C1_040_net_fail
+ C0_041_net_fail C1_041_net_fail
+ C0_042_net_fail C1_042_net_fail
+ C0_043_net_fail C1_043_net_fail
+ C0_044_net_fail C1_044_net_fail
+ C0_045_net_fail C1_045_net_fail
+ C0_046_net_fail C1_046_net_fail
+ C0_047_net_fail C1_047_net_fail
+ C0_048_net_fail C1_048_net_fail
+ C0_049_net_fail C1_049_net_fail
+ C0_050_net_fail C1_050_net_fail
+ C0_051_net_fail C1_051_net_fail
+ C0_052_net_fail C1_052_net_fail
+ C0_053_net_fail C1_053_net_fail
+ C0_054_net_fail C1_054_net_fail
+ C0_055_net_fail C1_055_net_fail
+ C0_056_net_fail C1_056_net_fail
+ C0_057_net_fail C1_057_net_fail
+ C0_058_net_fail C1_058_net_fail
+ C0_059_net_fail C1_059_net_fail
+ C0_060_net_fail C1_060_net_fail
+ C0_061_net_fail C1_061_net_fail
+ C0_062_net_fail C1_062_net_fail
+ C0_063_net_fail C1_063_net_fail

C000_net_fail C0_000_net_fail C1_000_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=0.22221p P=2.91342u

C001_net_fail C0_001_net_fail C1_001_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=0.44442p P=5.38242u

C002_net_fail C0_002_net_fail C1_002_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=0.6666300000000001p P=7.85142u

C003_net_fail C0_003_net_fail C1_003_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=0.88884p P=10.320419999999999u

C004_net_fail C0_004_net_fail C1_004_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=0.44442p P=3.35784u

C005_net_fail C0_005_net_fail C1_005_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=0.88884p P=5.82684u

C006_net_fail C0_006_net_fail C1_006_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=1.3332600000000001p P=8.29584u

C007_net_fail C0_007_net_fail C1_007_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=1.77768p P=10.76484u

C008_net_fail C0_008_net_fail C1_008_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=0.6666300000000001p P=3.80226u

C009_net_fail C0_009_net_fail C1_009_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=1.3332600000000001p P=6.27126u

C010_net_fail C0_010_net_fail C1_010_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=1.99989p P=8.74026u

C011_net_fail C0_011_net_fail C1_011_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=2.6665200000000002p P=11.209259999999999u

C012_net_fail C0_012_net_fail C1_012_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=0.88884p P=4.24668u

C013_net_fail C0_013_net_fail C1_013_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=1.77768p P=6.71568u

C014_net_fail C0_014_net_fail C1_014_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=2.6665200000000002p P=9.18468u

C015_net_fail C0_015_net_fail C1_015_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=3.55536p P=11.65368u

C016_net_fail C0_016_net_fail C1_016_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=1.1110499999999999p P=14.5671u

C017_net_fail C0_017_net_fail C1_017_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=2.2220999999999997p P=26.9121u

C018_net_fail C0_018_net_fail C1_018_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=3.33315p P=39.2571u

C019_net_fail C0_019_net_fail C1_019_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=4.4441999999999995p P=51.60209999999999u

C020_net_fail C0_020_net_fail C1_020_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=2.2220999999999997p P=16.789199999999997u

C021_net_fail C0_021_net_fail C1_021_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=4.4441999999999995p P=29.1342u

C022_net_fail C0_022_net_fail C1_022_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=6.6663p P=41.4792u

C023_net_fail C0_023_net_fail C1_023_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=8.888399999999999p P=53.8242u

C024_net_fail C0_024_net_fail C1_024_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=3.33315p P=19.0113u

C025_net_fail C0_025_net_fail C1_025_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=6.6663p P=31.356299999999997u

C026_net_fail C0_026_net_fail C1_026_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=9.99945p P=43.701299999999996u

C027_net_fail C0_027_net_fail C1_027_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=13.3326p P=56.046299999999995u

C028_net_fail C0_028_net_fail C1_028_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=4.4441999999999995p P=21.2334u

C029_net_fail C0_029_net_fail C1_029_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=8.888399999999999p P=33.578399999999995u

C030_net_fail C0_030_net_fail C1_030_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=13.3326p P=45.9234u

C031_net_fail C0_031_net_fail C1_031_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=17.776799999999998p P=58.2684u

C032_net_fail C0_032_net_fail C1_032_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=1.99989p P=26.220779999999998u

C033_net_fail C0_033_net_fail C1_033_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=3.99978p P=48.44178u

C034_net_fail C0_034_net_fail C1_034_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=5.99967p P=70.66278u

C035_net_fail C0_035_net_fail C1_035_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=7.99956p P=92.88377999999999u

C036_net_fail C0_036_net_fail C1_036_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=3.99978p P=30.22056u

C037_net_fail C0_037_net_fail C1_037_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=7.99956p P=52.441559999999996u

C038_net_fail C0_038_net_fail C1_038_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=11.99934p P=74.66255999999998u

C039_net_fail C0_039_net_fail C1_039_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=15.99912p P=96.88356u

C040_net_fail C0_040_net_fail C1_040_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=5.99967p P=34.22034u

C041_net_fail C0_041_net_fail C1_041_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=11.99934p P=56.44134u

C042_net_fail C0_042_net_fail C1_042_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=17.99901p P=78.66234u

C043_net_fail C0_043_net_fail C1_043_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=23.99868p P=100.88333999999999u

C044_net_fail C0_044_net_fail C1_044_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=7.99956p P=38.22012u

C045_net_fail C0_045_net_fail C1_045_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=15.99912p P=60.44112u

C046_net_fail C0_046_net_fail C1_046_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=23.99868p P=82.66211999999999u

C047_net_fail C0_047_net_fail C1_047_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=31.99824p P=104.88311999999999u

C048_net_fail C0_048_net_fail C1_048_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=2.88873p P=37.87446u

C049_net_fail C0_049_net_fail C1_049_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=5.77746p P=69.97146u

C050_net_fail C0_050_net_fail C1_050_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=8.666189999999999p P=102.06846u

C051_net_fail C0_051_net_fail C1_051_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=11.55492p P=134.16546u

C052_net_fail C0_052_net_fail C1_052_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=5.77746p P=43.65192u

C053_net_fail C0_053_net_fail C1_053_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=11.55492p P=75.74892u

C054_net_fail C0_054_net_fail C1_054_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=17.332379999999997p P=107.84591999999999u

C055_net_fail C0_055_net_fail C1_055_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=23.10984p P=139.94292u

C056_net_fail C0_056_net_fail C1_056_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=8.666189999999999p P=49.429379999999995u

C057_net_fail C0_057_net_fail C1_057_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=17.332379999999997p P=81.52638u

C058_net_fail C0_058_net_fail C1_058_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=25.998569999999997p P=113.62338u

C059_net_fail C0_059_net_fail C1_059_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=34.664759999999994p P=145.72038u

C060_net_fail C0_060_net_fail C1_060_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=11.55492p P=55.20683999999999u

C061_net_fail C0_061_net_fail C1_061_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=23.10984p P=87.30384u

C062_net_fail C0_062_net_fail C1_062_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=34.664759999999994p P=119.40083999999999u

C063_net_fail C0_063_net_fail C1_063_net_fail SUBSTRATE sky130_fd_pr__cap_var_hvt A=46.21968p P=151.49784u

.ENDS