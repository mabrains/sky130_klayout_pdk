*** LS Include files.

.include ./ls_cdl/sky130_fd_sc_ls__a2111o_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a2111o_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a2111o_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a2111oi_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a2111oi_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a2111oi_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a211o_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a211o_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a211o_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a211oi_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a211oi_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a211oi_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a21bo_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a21bo_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a21bo_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a21boi_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a21boi_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a21boi_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a21o_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a21o_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a21o_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a21oi_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a21oi_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a21oi_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a221o_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a221o_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a221o_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a221oi_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a221oi_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a221oi_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a222o_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a222o_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a222oi_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a222oi_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a22o_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a22o_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a22o_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a22oi_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a22oi_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a22oi_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a2bb2o_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a2bb2o_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a2bb2o_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a2bb2oi_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a2bb2oi_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a2bb2oi_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a311o_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a311o_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a311o_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a311oi_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a311oi_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a311oi_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a31o_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a31o_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a31o_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a31oi_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a31oi_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a31oi_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a32o_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a32o_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a32o_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a32oi_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a32oi_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a32oi_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a41o_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a41o_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a41o_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a41oi_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a41oi_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__a41oi_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and2_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and2_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and2_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and2b_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and2b_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and2b_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and3_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and3_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and3_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and3b_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and3b_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and3b_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and4_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and4_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and4_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and4b_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and4b_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and4b_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and4bb_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and4bb_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__and4bb_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__buf_16.cdl
.include ./ls_cdl/sky130_fd_sc_ls__buf_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__buf_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__buf_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__buf_8.cdl
.include ./ls_cdl/sky130_fd_sc_ls__bufbuf_16.cdl
.include ./ls_cdl/sky130_fd_sc_ls__bufbuf_8.cdl
.include ./ls_cdl/sky130_fd_sc_ls__bufinv_16.cdl
.include ./ls_cdl/sky130_fd_sc_ls__bufinv_8.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkbuf_16.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkbuf_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkbuf_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkbuf_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkbuf_8.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkdlyinv3sd1_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkdlyinv3sd2_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkdlyinv3sd3_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkdlyinv5sd1_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkdlyinv5sd2_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkdlyinv5sd3_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkinv_16.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkinv_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkinv_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkinv_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__clkinv_8.cdl
.include ./ls_cdl/sky130_fd_sc_ls__decap_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__decap_8.cdl
.include ./ls_cdl/sky130_fd_sc_ls__decaphe_18.cdl
.include ./ls_cdl/sky130_fd_sc_ls__decaphe_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__decaphe_3.cdl
.include ./ls_cdl/sky130_fd_sc_ls__decaphe_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__decaphe_6.cdl
.include ./ls_cdl/sky130_fd_sc_ls__decaphe_8.cdl
.include ./ls_cdl/sky130_fd_sc_ls__decaphetap_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfbbn_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfbbn_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfbbp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfrbp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfrbp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfrtn_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfrtp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfrtp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfrtp_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfsbp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfsbp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfstp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfstp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfstp_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfxbp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfxbp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfxtp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfxtp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dfxtp_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlclkp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlclkp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlclkp_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlrbn_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlrbn_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlrbp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlrbp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlrtn_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlrtn_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlrtn_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlrtp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlrtp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlrtp_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlxbn_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlxbn_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlxbp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlxtn_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlxtn_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlxtn_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlxtp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlygate4sd1_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlygate4sd2_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlygate4sd3_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlymetal6s2s_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlymetal6s4s_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__dlymetal6s6s_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__ebufn_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__ebufn_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__ebufn_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__ebufn_8.cdl
.include ./ls_cdl/sky130_fd_sc_ls__edfxbp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__edfxtp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__einvn_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__einvn_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__einvn_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__einvn_8.cdl
.include ./ls_cdl/sky130_fd_sc_ls__einvp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__einvp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__einvp_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__einvp_8.cdl
.include ./ls_cdl/sky130_fd_sc_ls__fa_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__fa_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__fa_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__fah_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__fah_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__fah_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__fahcin_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__fahcon_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__ha_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__ha_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__ha_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__inv_16.cdl
.include ./ls_cdl/sky130_fd_sc_ls__inv_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__inv_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__inv_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__inv_8.cdl
.include ./ls_cdl/sky130_fd_sc_ls__maj3_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__maj3_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__maj3_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__mux2_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__mux2_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__mux2_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__mux2i_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__mux2i_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__mux2i_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__mux4_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__mux4_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__mux4_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand2_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand2_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand2_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand2_8.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand2b_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand2b_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand2b_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand3_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand3_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand3_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand3b_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand3b_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand3b_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand4_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand4_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand4_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand4b_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand4b_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand4b_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand4bb_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand4bb_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nand4bb_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor2_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor2_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor2_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor2_8.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor2b_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor2b_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor2b_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor3_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor3_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor3_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor3b_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor3b_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor3b_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor4_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor4_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor4_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor4b_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor4b_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor4b_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor4bb_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor4bb_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__nor4bb_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o2111a_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o2111a_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o2111a_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o2111ai_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o2111ai_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o2111ai_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o211a_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o211a_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o211a_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o211ai_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o211ai_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o211ai_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o21a_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o21a_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o21a_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o21ai_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o21ai_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o21ai_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o21ba_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o21ba_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o21ba_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o21bai_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o21bai_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o21bai_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o221a_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o221a_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o221a_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o221ai_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o221ai_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o221ai_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o22a_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o22a_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o22a_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o22ai_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o22ai_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o22ai_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o2bb2a_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o2bb2a_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o2bb2a_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o2bb2ai_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o2bb2ai_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o2bb2ai_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o311a_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o311a_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o311a_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o311ai_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o311ai_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o311ai_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o31a_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o31a_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o31a_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o31ai_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o31ai_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o31ai_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o32a_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o32a_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o32a_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o32ai_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o32ai_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o32ai_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o41a_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o41a_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o41a_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o41ai_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o41ai_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__o41ai_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or2_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or2_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or2_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or2b_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or2b_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or2b_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or3_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or3_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or3_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or3b_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or3b_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or3b_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or4_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or4_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or4_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or4b_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or4b_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or4b_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or4bb_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or4bb_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__or4bb_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfbbn_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfbbn_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfbbp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfrbp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfrbp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfrtn_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfrtp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfrtp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfrtp_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfsbp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfsbp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfstp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfstp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfstp_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfxbp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfxbp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfxtp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfxtp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdfxtp_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdlclkp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdlclkp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sdlclkp_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sedfxbp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sedfxbp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sedfxtp_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sedfxtp_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__sedfxtp_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__xnor2_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__xnor2_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__xnor2_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__xnor3_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__xnor3_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__xnor3_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__xor2_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__xor2_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__xor2_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__xor3_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__xor3_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__xor3_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__conb_1.cdl
.include ./ls_cdl/sky130_fd_sc_ls__diode_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__fill_diode_2.cdl
.include ./ls_cdl/sky130_fd_sc_ls__fill_diode_4.cdl
.include ./ls_cdl/sky130_fd_sc_ls__fill_diode_8.cdl
