 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT diode 
+ D0_000 D1_000
+ D0_031 D1_031
+ D0_063 D1_063
+ D0_000 D1_000
+ D0_031 D1_031
+ D0_063 D1_063
+ D0_000 D1_000
+ D0_031 D1_031
+ D0_063 D1_063
+ D0_000 D1_000
+ D0_031 D1_031
+ D0_063 D1_063
+ D0_000 D1_000
+ D0_031 D1_031
+ D0_063 D1_063
+ D0_000 D1_000
+ D0_031 D1_031
+ D0_063 D1_063
+ D0_000 D1_000
+ D0_031 D1_031
+ D0_063 D1_063
+ D0_000 D1_000
+ D0_031 D1_031
+ D0_063 D1_063
+ D0 D1


D000 D0_000 D1_000 sky130_fd_pr__diode_pd2nw_05v5 AREA=0.2025 PJ=1.8

D031 D0_031 D1_031 sky130_fd_pr__diode_pd2nw_05v5 AREA=6.48 PJ=10.8

D063 D0_063 D1_063 sky130_fd_pr__diode_pd2nw_05v5 AREA=12.96 PJ=14.4

D000 D0_000 D1_000 sky130_fd_pr__diode_pd2nw_05v5_hvt AREA=0.2025 PJ=1.8

D031 D0_031 D1_031 sky130_fd_pr__diode_pd2nw_05v5_hvt AREA=6.48 PJ=10.8

D063 D0_063 D1_063 sky130_fd_pr__diode_pd2nw_05v5_hvt AREA=12.96 PJ=14.4

D000 D0_000 D1_000 sky130_fd_pr__diode_pd2nw_05v5_lvt AREA=0.2025 PJ=1.8

D031 D0_031 D1_031 sky130_fd_pr__diode_pd2nw_05v5_lvt AREA=6.48 PJ=10.8

D063 D0_063 D1_063 sky130_fd_pr__diode_pd2nw_05v5_lvt AREA=12.96 PJ=14.4

D000 D0_000 D1_000 sky130_fd_pr__diode_pd2nw_11v0 AREA=0.2025 PJ=1.8

D031 D0_031 D1_031 sky130_fd_pr__diode_pd2nw_11v0 AREA=6.48 PJ=10.8

D063 D0_063 D1_063 sky130_fd_pr__diode_pd2nw_11v0 AREA=12.96 PJ=14.4

D000 D0_000 D1_000 sky130_fd_pr__diode_pw2nd_05v5 AREA=0.2025 PJ=1.8

D031 D0_031 D1_031 sky130_fd_pr__diode_pw2nd_05v5 AREA=6.48 PJ=10.8

D063 D0_063 D1_063 sky130_fd_pr__diode_pw2nd_05v5 AREA=12.96 PJ=14.4

D000 D0_000 D1_000 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=0.2025 PJ=1.8

D031 D0_031 D1_031 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=6.48 PJ=10.8

D063 D0_063 D1_063 sky130_fd_pr__diode_pw2nd_05v5_lvt AREA=12.96 PJ=14.4

D000 D0_000 D1_000 sky130_fd_pr__diode_pw2nd_05v5_nvt AREA=0.2025 PJ=1.8

D031 D0_031 D1_031 sky130_fd_pr__diode_pw2nd_05v5_nvt AREA=6.48 PJ=10.8

D063 D0_063 D1_063 sky130_fd_pr__diode_pw2nd_05v5_nvt AREA=12.96 PJ=14.4

D000 D0_000 D1_000 sky130_fd_pr__diode_pw2nd_11v0 AREA=0.2025 PJ=1.8

D031 D0_031 D1_031 sky130_fd_pr__diode_pw2nd_11v0 AREA=6.48 PJ=10.8

D063 D0_063 D1_063 sky130_fd_pr__diode_pw2nd_11v0 AREA=12.96 PJ=14.4

Dx D0 D1 sky130_fd_pr__photodiode

.ENDS