* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_lp__dlybuf4s50kapwr_2 A KAPWR VGND VNB VPB VPWR X
*.PININFO A:I KAPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIP1 X Ab KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.26U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMIP0 net56 A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI10 net52 net56 KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI12 Ab net52 KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI7 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.42U l=0.15U mult=1 sa=0.265 sb=0.265
+ sd=0.28 area=0.063 perim=1.14
MMIN0 net56 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI9 net52 net56 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=1.0U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI11 Ab net52 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=1.0U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
.ENDS sky130_fd_sc_lp__dlybuf4s50kapwr_2
