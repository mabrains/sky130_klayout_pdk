*** LP Include files.

.include ./lp_cdl/sky130_fd_sc_lp__a2111o_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2111o_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2111o_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2111o_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2111oi_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2111oi_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2111oi_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2111oi_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2111oi_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2111oi_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2111o_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2111o_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a211o_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a211o_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a211o_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a211o_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a211oi_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a211oi_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a211oi_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a211oi_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a211oi_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a211oi_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a211o_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a211o_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21bo_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21bo_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21bo_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21bo_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21boi_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21boi_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21boi_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21boi_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21boi_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21boi_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21bo_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21bo_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21o_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21o_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21o_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21o_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21oi_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21oi_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21oi_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21oi_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21oi_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21oi_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21o_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a21o_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a221o_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a221o_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a221o_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a221o_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a221oi_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a221oi_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a221oi_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a221oi_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a221oi_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a221oi_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a221o_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a221o_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a22o_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a22o_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a22o_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a22o_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a22oi_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a22oi_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a22oi_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a22oi_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a22oi_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a22oi_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a22o_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a22o_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2bb2o_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2bb2o_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2bb2o_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2bb2o_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2bb2oi_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2bb2oi_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2bb2oi_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2bb2oi_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2bb2oi_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2bb2oi_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2bb2o_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a2bb2o_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a311o_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a311o_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a311o_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a311o_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a311oi_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a311oi_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a311oi_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a311oi_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a311oi_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a311oi_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a311o_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a311o_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a31o_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a31o_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a31o_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a31o_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a31oi_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a31oi_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a31oi_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a31oi_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a31oi_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a31oi_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a31o_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a31o_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a32o_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a32o_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a32o_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a32o_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a32oi_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a32oi_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a32oi_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a32oi_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a32oi_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a32oi_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a32o_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a32o_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a41o_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a41o_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a41o_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a41o_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a41oi_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a41oi_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a41oi_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a41oi_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a41oi_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a41oi_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a41o_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__a41o_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and2_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and2_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and2_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and2_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and2b_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and2b_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and2b_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and2b_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and2b_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and2_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and2_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and2_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and3_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and3_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and3_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and3_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and3b_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and3b_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and3b_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and3b_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and3b_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and3_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and3_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4b_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4b_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4b_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4bb_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4bb_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4bb_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4bb_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4bb_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4b_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4b_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__and4_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__buf_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__buf_16.cdl
.include ./lp_cdl/sky130_fd_sc_lp__buf_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__buf_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__buf_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__buf_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__bufbuf_16.cdl
.include ./lp_cdl/sky130_fd_sc_lp__bufbuf_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__bufinv_16.cdl
.include ./lp_cdl/sky130_fd_sc_lp__bufinv_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__bufkapwr_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__bufkapwr_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__bufkapwr_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__bufkapwr_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__buflp_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__buflp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__buflp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__buflp_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__buflp_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__buf_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__buflp_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__buf_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__busdriver_20.cdl
.include ./lp_cdl/sky130_fd_sc_lp__busdriver2_20.cdl
.include ./lp_cdl/sky130_fd_sc_lp__busdrivernovlp_20.cdl
.include ./lp_cdl/sky130_fd_sc_lp__busdrivernovlp2_20.cdl
.include ./lp_cdl/sky130_fd_sc_lp__busdrivernovlpsleep_20.cdl
.include ./lp_cdl/sky130_fd_sc_lp__bushold0_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__bushold_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__busreceiver_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__busreceiver_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__busreceiver_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkbuf_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkbuf_16.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkbuf_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkbuf_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkbuf_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkbuf_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkbuf_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkdlybuf4s15_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkdlybuf4s15_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkdlybuf4s18_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkdlybuf4s18_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkdlybuf4s25_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkdlybuf4s25_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkdlybuf4s50_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkdlybuf4s50_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkinv_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkinv_16.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkinv_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkinv_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkinv_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkinv_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkinv_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkinvlp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkinv_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__conb_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__conb_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__decap_12.cdl
.include ./lp_cdl/sky130_fd_sc_lp__decap_3.cdl
.include ./lp_cdl/sky130_fd_sc_lp__decap_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__decap_6.cdl
.include ./lp_cdl/sky130_fd_sc_lp__decap_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__decapkapwr_12.cdl
.include ./lp_cdl/sky130_fd_sc_lp__decapkapwr_3.cdl
.include ./lp_cdl/sky130_fd_sc_lp__decapkapwr_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__decapkapwr_6.cdl
.include ./lp_cdl/sky130_fd_sc_lp__decapkapwr_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfbbn_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfbbn_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfbbp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfrbp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfrbp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfrbp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfrtn_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfrtp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfrtp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfrtp_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfsbp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfsbp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfsbp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfstp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfstp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfstp_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfstp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfxbp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfxbp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfxbp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfxtp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfxtp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfxtp_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dfxtp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlclkp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlclkp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlclkp_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlclkp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlrbn_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlrbn_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlrbn_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlrbp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlrbp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlrbp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlrtn_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlrtn_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlrtn_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlrtn_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlrtp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlrtp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlrtp_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlrtp_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlrtp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlxbn_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlxbn_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlxbp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlxbp_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlxbp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlxtn_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlxtn_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlxtn_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlxtp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlxtp_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlxtp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlybuf4s15kapwr_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlybuf4s15kapwr_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlybuf4s18kapwr_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlybuf4s18kapwr_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlybuf4s25kapwr_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlybuf4s25kapwr_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlybuf4s50kapwr_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlybuf4s50kapwr_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlygate4s15_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlygate4s18_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlygate4s50_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlymetal6s2s_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlymetal6s4s_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__dlymetal6s6s_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__ebufn_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__ebufn_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__ebufn_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__ebufn_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__ebufn_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__ebufn_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__edfxbp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__einvn_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__einvn_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__einvn_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__einvn_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__einvn_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__einvn_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__einvn_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__einvp_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__einvp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__einvp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__einvp_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__einvp_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__einvp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__einvp_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__fa_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__fa_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__fa_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__fa_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__fah_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__fahcin_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__fahcon_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__fa_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__fa_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__ha_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__ha_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__ha_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__ha_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__ha_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__ha_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__inputiso0n_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__inputiso0p_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__inputiso1n_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__inputiso1p_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__inputisolatch_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__inv_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__inv_16.cdl
.include ./lp_cdl/sky130_fd_sc_lp__inv_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__inv_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__inv_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__inv_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__invkapwr_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__invkapwr_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__invkapwr_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__invkapwr_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__invlp_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__invlp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__invlp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__invlp_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__invlp_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__inv_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__invlp_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__inv_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__iso0n_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__iso0n_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__iso0p_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__iso0p_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__iso1n_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__iso1n_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__iso1p_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__iso1p_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__isobufsrc_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__isobufsrc_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__isobufsrc_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__isolatch_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__lsbufiso0p_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__lsbufiso1p_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__lsbuf_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__maj3_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__maj3_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__maj3_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__maj3_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__maj3_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__maj3_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux2_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux2_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux2_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux2_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux2_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux2i_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux2i_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux2i_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux2i_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux2i_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux2i_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux2i_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux2_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux2_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux2_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux4_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux4_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux4_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux4_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux4_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__mux4_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand2_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand2_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand2_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand2_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand2_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand2b_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand2b_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand2b_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand2b_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand2b_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand2_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand2_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand2_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand3_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand3_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand3_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand3_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand3b_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand3b_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand3b_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand3b_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand3b_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand3_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand3_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4b_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4b_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4b_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4bb_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4bb_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4bb_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4bb_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4bb_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4b_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4b_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nand4_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor2_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor2_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor2_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor2_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor2_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor2b_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor2b_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor2b_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor2b_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor2b_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor2_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor2_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor2_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor3_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor3_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor3_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor3_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor3b_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor3b_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor3b_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor3b_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor3b_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor3_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor3_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4b_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4b_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4b_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4bb_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4bb_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4bb_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4bb_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4bb_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4b_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4b_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__nor4_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2111a_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2111a_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2111a_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2111a_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2111ai_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2111ai_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2111ai_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2111ai_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2111ai_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2111ai_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2111a_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2111a_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o211a_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o211a_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o211a_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o211a_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o211ai_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o211ai_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o211ai_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o211ai_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o211ai_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o211ai_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o211a_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o211a_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21a_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21a_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21a_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21a_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21ai_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21ai_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21ai_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21ai_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21ai_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21ai_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21a_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21a_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21ba_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21ba_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21ba_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21ba_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21bai_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21bai_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21bai_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21bai_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21bai_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21bai_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21ba_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o21ba_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o221a_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o221a_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o221a_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o221a_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o221ai_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o221ai_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o221ai_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o221ai_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o221ai_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o221ai_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o221a_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o221a_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o22a_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o22a_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o22a_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o22a_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o22ai_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o22ai_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o22ai_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o22ai_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o22ai_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o22ai_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o22a_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o22a_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2bb2a_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2bb2a_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2bb2a_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2bb2a_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2bb2ai_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2bb2ai_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2bb2ai_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2bb2ai_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2bb2ai_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2bb2ai_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2bb2a_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o2bb2a_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o311a_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o311a_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o311a_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o311a_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o311ai_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o311ai_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o311ai_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o311ai_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o311ai_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o311ai_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o311a_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o311a_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o31a_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o31a_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o31a_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o31a_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o31ai_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o31ai_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o31ai_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o31ai_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o31ai_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o31ai_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o31a_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o31a_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o32a_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o32a_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o32a_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o32a_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o32ai_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o32ai_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o32ai_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o32ai_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o32ai_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o32ai_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o32a_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o32a_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o41a_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o41a_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o41a_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o41a_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o41ai_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o41ai_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o41ai_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o41ai_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o41ai_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o41ai_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o41a_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__o41a_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or2_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or2_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or2_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or2_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or2b_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or2b_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or2b_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or2b_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or2b_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or2_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or2_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or2_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or3_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or3_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or3_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or3_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or3b_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or3b_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or3b_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or3b_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or3b_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or3_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or3_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4b_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4b_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4b_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4bb_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4bb_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4bb_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4bb_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4bb_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4b_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4b_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__or4_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfbbn_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfbbn_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfbbp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfrbp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfrbp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfrbp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfrtn_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfrtp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfrtp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfrtp_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfrtp_lp2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfrtp_ov2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfsbp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfsbp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfsbp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfstp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfstp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfstp_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfstp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfxbp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfxbp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfxbp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfxtp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfxtp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfxtp_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdfxtp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdlclkp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdlclkp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdlclkp_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sdlclkp_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sleep_pargate_plv_14.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sleep_pargate_plv_21.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sleep_pargate_plv_28.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sleep_pargate_plv_7.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sleep_sergate_plv_14.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sleep_sergate_plv_21.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sleep_sergate_plv_28.cdl
.include ./lp_cdl/sky130_fd_sc_lp__srdlrtp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__srdlstp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__srdlxtp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sregrbp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__sregsbp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__srsdfrtn_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__srsdfrtp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__srsdfstp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__srsdfxtp_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xnor2_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xnor2_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xnor2_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xnor2_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xnor2_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xnor2_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xnor3_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xnor3_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xor2_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xor2_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xor2_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xor2_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xor2_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xor2_m.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xor3_1.cdl
.include ./lp_cdl/sky130_fd_sc_lp__xor3_lp.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkbuflp_16.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkbuflp_2.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkbuflp_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkbuflp_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkinvlp_16.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkinvlp_4.cdl
.include ./lp_cdl/sky130_fd_sc_lp__clkinvlp_8.cdl
.include ./lp_cdl/sky130_fd_sc_lp__diode_0.cdl
.include ./lp_cdl/sky130_fd_sc_lp__diode_1.cdl
