* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hdll__xor2_1 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMNnor0 inor A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0U l=0.18U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0U l=0.18U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0U l=0.18U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0U l=0.18U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0U l=0.18U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_hdll__xor2_1
