 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__res_xhigh_po_5p73
+ R0_0 R1_0
+ R0_1 R1_1
+ R0_2 R1_2
+ R0_3 R1_3
+ R0_4 R1_4
+ R0_5 R1_5
+ R0_6 R1_6
+ R0_7 R1_7
+ R0_8 R1_8
+ R0_9 R1_9
+ R0_10 R1_10
+ R0_11 R1_11
+ R0_12 R1_12
+ R0_13 R1_13
+ R0_14 R1_14
+ R0_15 R1_15
+ R0_16 R1_16
+ R0_17 R1_17
+ R0_18 R1_18
+ R0_19 R1_19
+ R0_20 R1_20
+ R0_21 R1_21
+ R0_22 R1_22
+ R0_23 R1_23
+ R0_24 R1_24
+ R0_25 R1_25
+ R0_26 R1_26
+ R0_27 R1_27
+ R0_28 R1_28
+ R0_29 R1_29
+ R0_30 R1_30
+ R0_31 R1_31
+ R0_32 R1_32
+ R0_33 R1_33
+ R0_34 R1_34
+ R0_35 R1_35
+ R0_36 R1_36
+ R0_37 R1_37
+ R0_38 R1_38
+ R0_39 R1_39
+ R0_40 R1_40
+ R0_41 R1_41
+ R0_42 R1_42
+ R0_43 R1_43
+ R0_44 R1_44
+ R0_45 R1_45
+ R0_46 R1_46
+ R0_47 R1_47
+ R0_48 R1_48
+ R0_49 R1_49
+ R0_50 R1_50
+ R0_51 R1_51
+ R0_52 R1_52
+ R0_53 R1_53
+ R0_54 R1_54
+ R0_55 R1_55
+ R0_56 R1_56
+ R0_57 R1_57
+ R0_58 R1_58
+ R0_59 R1_59
+ R0_60 R1_60
+ R0_61 R1_61
+ R0_62 R1_62
+ R0_63 R1_63

R0 R0_0 R1_0 sky130_fd_pr__res_xhigh_po_5p73 l=6.23 w=5.73

R1 R0_1 R1_1 sky130_fd_pr__res_xhigh_po_5p73 l=12.46 w=5.73

R2 R0_2 R1_2 sky130_fd_pr__res_xhigh_po_5p73 l=18.69 w=5.73

R3 R0_3 R1_3 sky130_fd_pr__res_xhigh_po_5p73 l=24.92 w=5.73

R4 R0_4 R1_4 sky130_fd_pr__res_xhigh_po_5p73 l=31.15 w=5.73

R5 R0_5 R1_5 sky130_fd_pr__res_xhigh_po_5p73 l=37.38 w=5.73

R6 R0_6 R1_6 sky130_fd_pr__res_xhigh_po_5p73 l=43.61 w=5.73

R7 R0_7 R1_7 sky130_fd_pr__res_xhigh_po_5p73 l=49.84 w=5.73

R8 R0_8 R1_8 sky130_fd_pr__res_xhigh_po_5p73 l=12.46 w=5.73

R9 R0_9 R1_9 sky130_fd_pr__res_xhigh_po_5p73 l=24.92 w=5.73

R10 R0_10 R1_10 sky130_fd_pr__res_xhigh_po_5p73 l=37.38 w=5.73

R11 R0_11 R1_11 sky130_fd_pr__res_xhigh_po_5p73 l=49.84 w=5.73

R12 R0_12 R1_12 sky130_fd_pr__res_xhigh_po_5p73 l=62.3 w=5.73

R13 R0_13 R1_13 sky130_fd_pr__res_xhigh_po_5p73 l=74.76 w=5.73

R14 R0_14 R1_14 sky130_fd_pr__res_xhigh_po_5p73 l=87.22 w=5.73

R15 R0_15 R1_15 sky130_fd_pr__res_xhigh_po_5p73 l=99.68 w=5.73

R16 R0_16 R1_16 sky130_fd_pr__res_xhigh_po_5p73 l=18.69 w=5.73

R17 R0_17 R1_17 sky130_fd_pr__res_xhigh_po_5p73 l=37.38 w=5.73

R18 R0_18 R1_18 sky130_fd_pr__res_xhigh_po_5p73 l=56.07 w=5.73

R19 R0_19 R1_19 sky130_fd_pr__res_xhigh_po_5p73 l=74.76 w=5.73

R20 R0_20 R1_20 sky130_fd_pr__res_xhigh_po_5p73 l=93.45 w=5.73

R21 R0_21 R1_21 sky130_fd_pr__res_xhigh_po_5p73 l=112.14 w=5.73

R22 R0_22 R1_22 sky130_fd_pr__res_xhigh_po_5p73 l=130.83 w=5.73

R23 R0_23 R1_23 sky130_fd_pr__res_xhigh_po_5p73 l=149.52 w=5.73

R24 R0_24 R1_24 sky130_fd_pr__res_xhigh_po_5p73 l=24.92 w=5.73

R25 R0_25 R1_25 sky130_fd_pr__res_xhigh_po_5p73 l=49.84 w=5.73

R26 R0_26 R1_26 sky130_fd_pr__res_xhigh_po_5p73 l=74.76 w=5.73

R27 R0_27 R1_27 sky130_fd_pr__res_xhigh_po_5p73 l=99.68 w=5.73

R28 R0_28 R1_28 sky130_fd_pr__res_xhigh_po_5p73 l=124.6 w=5.73

R29 R0_29 R1_29 sky130_fd_pr__res_xhigh_po_5p73 l=149.52 w=5.73

R30 R0_30 R1_30 sky130_fd_pr__res_xhigh_po_5p73 l=174.44 w=5.73

R31 R0_31 R1_31 sky130_fd_pr__res_xhigh_po_5p73 l=199.36 w=5.73

R32 R0_32 R1_32 sky130_fd_pr__res_xhigh_po_5p73 l=31.15 w=5.73

R33 R0_33 R1_33 sky130_fd_pr__res_xhigh_po_5p73 l=62.3 w=5.73

R34 R0_34 R1_34 sky130_fd_pr__res_xhigh_po_5p73 l=93.45 w=5.73

R35 R0_35 R1_35 sky130_fd_pr__res_xhigh_po_5p73 l=124.6 w=5.73

R36 R0_36 R1_36 sky130_fd_pr__res_xhigh_po_5p73 l=155.75 w=5.73

R37 R0_37 R1_37 sky130_fd_pr__res_xhigh_po_5p73 l=186.9 w=5.73

R38 R0_38 R1_38 sky130_fd_pr__res_xhigh_po_5p73 l=218.05 w=5.73

R39 R0_39 R1_39 sky130_fd_pr__res_xhigh_po_5p73 l=249.2 w=5.73

R40 R0_40 R1_40 sky130_fd_pr__res_xhigh_po_5p73 l=37.38 w=5.73

R41 R0_41 R1_41 sky130_fd_pr__res_xhigh_po_5p73 l=74.76 w=5.73

R42 R0_42 R1_42 sky130_fd_pr__res_xhigh_po_5p73 l=112.14 w=5.73

R43 R0_43 R1_43 sky130_fd_pr__res_xhigh_po_5p73 l=149.52 w=5.73

R44 R0_44 R1_44 sky130_fd_pr__res_xhigh_po_5p73 l=186.9 w=5.73

R45 R0_45 R1_45 sky130_fd_pr__res_xhigh_po_5p73 l=224.28 w=5.73

R46 R0_46 R1_46 sky130_fd_pr__res_xhigh_po_5p73 l=261.66 w=5.73

R47 R0_47 R1_47 sky130_fd_pr__res_xhigh_po_5p73 l=299.04 w=5.73

R48 R0_48 R1_48 sky130_fd_pr__res_xhigh_po_5p73 l=43.61 w=5.73

R49 R0_49 R1_49 sky130_fd_pr__res_xhigh_po_5p73 l=87.22 w=5.73

R50 R0_50 R1_50 sky130_fd_pr__res_xhigh_po_5p73 l=130.83 w=5.73

R51 R0_51 R1_51 sky130_fd_pr__res_xhigh_po_5p73 l=174.44 w=5.73

R52 R0_52 R1_52 sky130_fd_pr__res_xhigh_po_5p73 l=218.05 w=5.73

R53 R0_53 R1_53 sky130_fd_pr__res_xhigh_po_5p73 l=261.66 w=5.73

R54 R0_54 R1_54 sky130_fd_pr__res_xhigh_po_5p73 l=305.27 w=5.73

R55 R0_55 R1_55 sky130_fd_pr__res_xhigh_po_5p73 l=348.88 w=5.73

R56 R0_56 R1_56 sky130_fd_pr__res_xhigh_po_5p73 l=49.84 w=5.73

R57 R0_57 R1_57 sky130_fd_pr__res_xhigh_po_5p73 l=99.68 w=5.73

R58 R0_58 R1_58 sky130_fd_pr__res_xhigh_po_5p73 l=149.52 w=5.73

R59 R0_59 R1_59 sky130_fd_pr__res_xhigh_po_5p73 l=199.36 w=5.73

R60 R0_60 R1_60 sky130_fd_pr__res_xhigh_po_5p73 l=249.2 w=5.73

R61 R0_61 R1_61 sky130_fd_pr__res_xhigh_po_5p73 l=299.04 w=5.73

R62 R0_62 R1_62 sky130_fd_pr__res_xhigh_po_5p73 l=348.88 w=5.73

R63 R0_63 R1_63 sky130_fd_pr__res_xhigh_po_5p73 l=398.72 w=5.73

.ENDS