* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI120 db SCE n1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.525 perim=3.1
MI103 n1 SCD VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.525 perim=3.1
MI104 db sceb n0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.525 perim=3.1
MI98 n0 D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.525 perim=3.1
MI657 M0 clkpos net72 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI656 net72 M1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI49 sceb SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI646 Q S1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI648 db clkneg M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI642 S0 clkneg net48 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI641 net48 S1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI649 S1 S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI634 M1 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI101 db sceb p1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI94 db D p0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI659 M0 clkneg net100 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI50 sceb SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI644 S0 clkpos net119 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI643 net119 S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI658 net100 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI645 Q S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI651 db clkpos M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
.ENDS sky130_fd_sc_hvl__sdfxtp_1
