* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_ms__dfsbp_2 CLK D SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI36 net64 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8_lvt m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net79 VNB nfet_01v8_lvt m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net111 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net64 VNB nfet_01v8_lvt m=1 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net96 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net104 VNB nfet_01v8_lvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net104 S1 net96 VNB nfet_01v8_lvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net111 VNB nfet_01v8_lvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net79 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net188 S0 VGND VNB nfet_01v8_lvt m=1 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net188 VGND VNB nfet_01v8_lvt m=2 w=0.74U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 Q_N S0 VGND VNB nfet_01v8_lvt m=2 w=0.74U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8 m=1 w=0.42U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net135 VPB pfet_01v8 m=1 w=1.0U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net135 M0 VPWR VPB pfet_01v8 m=1 w=1.0U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12U l=0.18U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.42U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net160 M1 VPWR VPB pfet_01v8 m=1 w=0.42U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net160 VPB pfet_01v8 m=1 w=0.42U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net171 S1 VPWR VPB pfet_01v8 m=1 w=0.42U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net171 VPB pfet_01v8 m=1 w=0.42U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8 m=1 w=0.42U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8 m=1 w=0.42U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.42U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net188 S0 VPWR VPB pfet_01v8 m=1 w=1.0U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net188 VPWR VPB pfet_01v8 m=2 w=1.12U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N S0 VPWR VPB pfet_01v8 m=2 w=1.12U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_ms__dfsbp_2
