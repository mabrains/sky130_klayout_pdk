* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_lp__sdfsbp_lp CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
MI645 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI663 net196 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI660 Q net196 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI661 Q_N S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI662 net111 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI664 M0 clkneg net111 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI6 net103 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI669 S0 clkpos net103 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI38 S0 clkneg net91 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI37 net91 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265 sb=0.265
+ sd=0.28 area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.25U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI34 S0 clkpos net224 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI27 net252 S1 net184 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI647 S1 S0 net180 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI655 M0 clkpos net243 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI656 M1 M0 net239 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI654 net243 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI676 net232 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI677 net228 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI36 net224 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI26 S0 clkneg net252 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI651 Q_N S0 net232 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI46 clkpos clkneg net164 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI44 clkneg CLK net172 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI657 net239 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI652 net196 S0 net228 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI644 sceb SCE net176 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI675 net188 net196 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI25 net184 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI674 net180 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI673 net176 SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI672 net172 CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI653 Q net196 net188 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI671 net164 clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265 sb=0.265
+ sd=0.28 area=0.525 perim=3.1
MI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.525 perim=3.1
MI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.525 perim=3.1
MI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.525 perim=3.1
.ENDS sky130_fd_sc_lp__sdfsbp_lp
