 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT res 
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063
+ R0_000 R1_000
+ R0_031 R1_031
+ R0_063 R1_063


R000 R0_000 R1_000 sky130_fd_pr__res_generic_l1 l=2.1 w=0.42

R031 R0_031 R1_031 sky130_fd_pr__res_generic_l1 l=8.4 w=3.36

R063 R0_063 R1_063 sky130_fd_pr__res_generic_l1 l=16.8 w=3.36

R000 R0_000 R1_000 sky130_fd_pr__res_generic_m1 l=2.1 w=0.42

R031 R0_031 R1_031 sky130_fd_pr__res_generic_m1 l=8.4 w=3.36

R063 R0_063 R1_063 sky130_fd_pr__res_generic_m1 l=16.8 w=3.36

R000 R0_000 R1_000 sky130_fd_pr__res_generic_m2 l=2.1 w=0.42

R031 R0_031 R1_031 sky130_fd_pr__res_generic_m2 l=8.4 w=3.36

R063 R0_063 R1_063 sky130_fd_pr__res_generic_m2 l=16.8 w=3.36

R000 R0_000 R1_000 sky130_fd_pr__res_generic_m3 l=2.1 w=0.42

R031 R0_031 R1_031 sky130_fd_pr__res_generic_m3 l=8.4 w=3.36

R063 R0_063 R1_063 sky130_fd_pr__res_generic_m3 l=16.8 w=3.36

R000 R0_000 R1_000 sky130_fd_pr__res_generic_m4 l=2.1 w=0.42

R031 R0_031 R1_031 sky130_fd_pr__res_generic_m4 l=8.4 w=3.36

R063 R0_063 R1_063 sky130_fd_pr__res_generic_m4 l=16.8 w=3.36

R000 R0_000 R1_000 sky130_fd_pr__res_generic_m5 l=2.1 w=0.42

R031 R0_031 R1_031 sky130_fd_pr__res_generic_m5 l=8.4 w=3.36

R063 R0_063 R1_063 sky130_fd_pr__res_generic_m5 l=16.8 w=3.36

R000 R0_000 R1_000 sky130_fd_pr__res_generic_nd l=2.1 w=0.42

R031 R0_031 R1_031 sky130_fd_pr__res_generic_nd l=8.4 w=3.36

R063 R0_063 R1_063 sky130_fd_pr__res_generic_nd l=16.8 w=3.36

R000 R0_000 R1_000 sky130_fd_pr__res_generic_nd_hv l=2.1 w=0.42

R031 R0_031 R1_031 sky130_fd_pr__res_generic_nd_hv l=8.4 w=3.36

R063 R0_063 R1_063 sky130_fd_pr__res_generic_nd_hv l=16.8 w=3.36

R000 R0_000 R1_000 sky130_fd_pr__res_generic_pd l=2.1 w=0.42

R031 R0_031 R1_031 sky130_fd_pr__res_generic_pd l=8.4 w=3.36

R063 R0_063 R1_063 sky130_fd_pr__res_generic_pd l=16.8 w=3.36

R000 R0_000 R1_000 sky130_fd_pr__res_generic_pd_hv l=2.1 w=0.42

R031 R0_031 R1_031 sky130_fd_pr__res_generic_pd_hv l=8.4 w=3.36

R063 R0_063 R1_063 sky130_fd_pr__res_generic_pd_hv l=16.8 w=3.36

R000 R0_000 R1_000 sky130_fd_pr__res_generic_po l=1.65 w=0.33

R031 R0_031 R1_031 sky130_fd_pr__res_generic_po l=6.6 w=2.64

R063 R0_063 R1_063 sky130_fd_pr__res_generic_po l=13.2 w=2.64

R000 R0_000 R1_000 sky130_fd_pr__res_high_po_0p35 l=0.85 w=0.35

R031 R0_031 R1_031 sky130_fd_pr__res_high_po_0p35 l=27.2 w=0.35

R063 R0_063 R1_063 sky130_fd_pr__res_high_po_0p35 l=54.4 w=0.35

R000 R0_000 R1_000 sky130_fd_pr__res_high_po_0p69 l=1.19 w=0.69

R031 R0_031 R1_031 sky130_fd_pr__res_high_po_0p69 l=38.08 w=0.69

R063 R0_063 R1_063 sky130_fd_pr__res_high_po_0p69 l=76.16 w=0.69

R000 R0_000 R1_000 sky130_fd_pr__res_high_po_1p41 l=1.91 w=1.41

R031 R0_031 R1_031 sky130_fd_pr__res_high_po_1p41 l=61.12 w=1.41

R063 R0_063 R1_063 sky130_fd_pr__res_high_po_1p41 l=122.24 w=1.41

R000 R0_000 R1_000 sky130_fd_pr__res_high_po_2p85 l=3.35 w=2.85

R031 R0_031 R1_031 sky130_fd_pr__res_high_po_2p85 l=107.2 w=2.85

R063 R0_063 R1_063 sky130_fd_pr__res_high_po_2p85 l=214.4 w=2.85

R000 R0_000 R1_000 sky130_fd_pr__res_high_po_5p73 l=6.23 w=5.73

R031 R0_031 R1_031 sky130_fd_pr__res_high_po_5p73 l=199.36 w=5.73

R063 R0_063 R1_063 sky130_fd_pr__res_high_po_5p73 l=398.72 w=5.73

R000 R0_000 R1_000 sky130_fd_pr__res_iso_pw l=26.5 w=2.65

R031 R0_031 R1_031 sky130_fd_pr__res_iso_pw l=106.0 w=21.2

R063 R0_063 R1_063 sky130_fd_pr__res_iso_pw l=212.0 w=21.2

R000 R0_000 R1_000 sky130_fd_pr__res_xhigh_po_0p35 l=0.85 w=0.35

R031 R0_031 R1_031 sky130_fd_pr__res_xhigh_po_0p35 l=27.2 w=0.35

R063 R0_063 R1_063 sky130_fd_pr__res_xhigh_po_0p35 l=54.4 w=0.35

R000 R0_000 R1_000 sky130_fd_pr__res_xhigh_po_0p69 l=1.19 w=0.69

R031 R0_031 R1_031 sky130_fd_pr__res_xhigh_po_0p69 l=38.08 w=0.69

R063 R0_063 R1_063 sky130_fd_pr__res_xhigh_po_0p69 l=76.16 w=0.69

R000 R0_000 R1_000 sky130_fd_pr__res_xhigh_po_1p41 l=1.91 w=1.41

R031 R0_031 R1_031 sky130_fd_pr__res_xhigh_po_1p41 l=61.12 w=1.41

R063 R0_063 R1_063 sky130_fd_pr__res_xhigh_po_1p41 l=122.24 w=1.41

R000 R0_000 R1_000 sky130_fd_pr__res_xhigh_po_2p85 l=3.35 w=2.85

R031 R0_031 R1_031 sky130_fd_pr__res_xhigh_po_2p85 l=107.2 w=2.85

R063 R0_063 R1_063 sky130_fd_pr__res_xhigh_po_2p85 l=214.4 w=2.85

R000 R0_000 R1_000 sky130_fd_pr__res_xhigh_po_5p73 l=6.23 w=5.73

R031 R0_031 R1_031 sky130_fd_pr__res_xhigh_po_5p73 l=199.36 w=5.73

R063 R0_063 R1_063 sky130_fd_pr__res_xhigh_po_5p73 l=398.72 w=5.73

.ENDS