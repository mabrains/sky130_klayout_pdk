 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__res_xhigh_po_2p85
+ R0_000 R1_000 R0_000_net_fail R0_000_dim_fail R1_000_net_fail R1_000_dim_fail
+ R0_001 R1_001 R0_001_net_fail R0_001_dim_fail R1_001_net_fail R1_001_dim_fail
+ R0_002 R1_002 R0_002_net_fail R0_002_dim_fail R1_002_net_fail R1_002_dim_fail
+ R0_003 R1_003 R0_003_net_fail R0_003_dim_fail R1_003_net_fail R1_003_dim_fail
+ R0_004 R1_004 R0_004_net_fail R0_004_dim_fail R1_004_net_fail R1_004_dim_fail
+ R0_005 R1_005 R0_005_net_fail R0_005_dim_fail R1_005_net_fail R1_005_dim_fail
+ R0_006 R1_006 R0_006_net_fail R0_006_dim_fail R1_006_net_fail R1_006_dim_fail
+ R0_007 R1_007 R0_007_net_fail R0_007_dim_fail R1_007_net_fail R1_007_dim_fail
+ R0_008 R1_008 R0_008_net_fail R0_008_dim_fail R1_008_net_fail R1_008_dim_fail
+ R0_009 R1_009 R0_009_net_fail R0_009_dim_fail R1_009_net_fail R1_009_dim_fail
+ R0_010 R1_010 R0_010_net_fail R0_010_dim_fail R1_010_net_fail R1_010_dim_fail
+ R0_011 R1_011 R0_011_net_fail R0_011_dim_fail R1_011_net_fail R1_011_dim_fail
+ R0_012 R1_012 R0_012_net_fail R0_012_dim_fail R1_012_net_fail R1_012_dim_fail
+ R0_013 R1_013 R0_013_net_fail R0_013_dim_fail R1_013_net_fail R1_013_dim_fail
+ R0_014 R1_014 R0_014_net_fail R0_014_dim_fail R1_014_net_fail R1_014_dim_fail
+ R0_015 R1_015 R0_015_net_fail R0_015_dim_fail R1_015_net_fail R1_015_dim_fail
+ R0_016 R1_016 R0_016_net_fail R0_016_dim_fail R1_016_net_fail R1_016_dim_fail
+ R0_017 R1_017 R0_017_net_fail R0_017_dim_fail R1_017_net_fail R1_017_dim_fail
+ R0_018 R1_018 R0_018_net_fail R0_018_dim_fail R1_018_net_fail R1_018_dim_fail
+ R0_019 R1_019 R0_019_net_fail R0_019_dim_fail R1_019_net_fail R1_019_dim_fail
+ R0_020 R1_020 R0_020_net_fail R0_020_dim_fail R1_020_net_fail R1_020_dim_fail
+ R0_021 R1_021 R0_021_net_fail R0_021_dim_fail R1_021_net_fail R1_021_dim_fail
+ R0_022 R1_022 R0_022_net_fail R0_022_dim_fail R1_022_net_fail R1_022_dim_fail
+ R0_023 R1_023 R0_023_net_fail R0_023_dim_fail R1_023_net_fail R1_023_dim_fail
+ R0_024 R1_024 R0_024_net_fail R0_024_dim_fail R1_024_net_fail R1_024_dim_fail
+ R0_025 R1_025 R0_025_net_fail R0_025_dim_fail R1_025_net_fail R1_025_dim_fail
+ R0_026 R1_026 R0_026_net_fail R0_026_dim_fail R1_026_net_fail R1_026_dim_fail
+ R0_027 R1_027 R0_027_net_fail R0_027_dim_fail R1_027_net_fail R1_027_dim_fail
+ R0_028 R1_028 R0_028_net_fail R0_028_dim_fail R1_028_net_fail R1_028_dim_fail
+ R0_029 R1_029 R0_029_net_fail R0_029_dim_fail R1_029_net_fail R1_029_dim_fail
+ R0_030 R1_030 R0_030_net_fail R0_030_dim_fail R1_030_net_fail R1_030_dim_fail
+ R0_031 R1_031 R0_031_net_fail R0_031_dim_fail R1_031_net_fail R1_031_dim_fail
+ R0_032 R1_032 R0_032_net_fail R0_032_dim_fail R1_032_net_fail R1_032_dim_fail
+ R0_033 R1_033 R0_033_net_fail R0_033_dim_fail R1_033_net_fail R1_033_dim_fail
+ R0_034 R1_034 R0_034_net_fail R0_034_dim_fail R1_034_net_fail R1_034_dim_fail
+ R0_035 R1_035 R0_035_net_fail R0_035_dim_fail R1_035_net_fail R1_035_dim_fail
+ R0_036 R1_036 R0_036_net_fail R0_036_dim_fail R1_036_net_fail R1_036_dim_fail
+ R0_037 R1_037 R0_037_net_fail R0_037_dim_fail R1_037_net_fail R1_037_dim_fail
+ R0_038 R1_038 R0_038_net_fail R0_038_dim_fail R1_038_net_fail R1_038_dim_fail
+ R0_039 R1_039 R0_039_net_fail R0_039_dim_fail R1_039_net_fail R1_039_dim_fail
+ R0_040 R1_040 R0_040_net_fail R0_040_dim_fail R1_040_net_fail R1_040_dim_fail
+ R0_041 R1_041 R0_041_net_fail R0_041_dim_fail R1_041_net_fail R1_041_dim_fail
+ R0_042 R1_042 R0_042_net_fail R0_042_dim_fail R1_042_net_fail R1_042_dim_fail
+ R0_043 R1_043 R0_043_net_fail R0_043_dim_fail R1_043_net_fail R1_043_dim_fail
+ R0_044 R1_044 R0_044_net_fail R0_044_dim_fail R1_044_net_fail R1_044_dim_fail
+ R0_045 R1_045 R0_045_net_fail R0_045_dim_fail R1_045_net_fail R1_045_dim_fail
+ R0_046 R1_046 R0_046_net_fail R0_046_dim_fail R1_046_net_fail R1_046_dim_fail
+ R0_047 R1_047 R0_047_net_fail R0_047_dim_fail R1_047_net_fail R1_047_dim_fail
+ R0_048 R1_048 R0_048_net_fail R0_048_dim_fail R1_048_net_fail R1_048_dim_fail
+ R0_049 R1_049 R0_049_net_fail R0_049_dim_fail R1_049_net_fail R1_049_dim_fail
+ R0_050 R1_050 R0_050_net_fail R0_050_dim_fail R1_050_net_fail R1_050_dim_fail
+ R0_051 R1_051 R0_051_net_fail R0_051_dim_fail R1_051_net_fail R1_051_dim_fail
+ R0_052 R1_052 R0_052_net_fail R0_052_dim_fail R1_052_net_fail R1_052_dim_fail
+ R0_053 R1_053 R0_053_net_fail R0_053_dim_fail R1_053_net_fail R1_053_dim_fail
+ R0_054 R1_054 R0_054_net_fail R0_054_dim_fail R1_054_net_fail R1_054_dim_fail
+ R0_055 R1_055 R0_055_net_fail R0_055_dim_fail R1_055_net_fail R1_055_dim_fail
+ R0_056 R1_056 R0_056_net_fail R0_056_dim_fail R1_056_net_fail R1_056_dim_fail
+ R0_057 R1_057 R0_057_net_fail R0_057_dim_fail R1_057_net_fail R1_057_dim_fail
+ R0_058 R1_058 R0_058_net_fail R0_058_dim_fail R1_058_net_fail R1_058_dim_fail
+ R0_059 R1_059 R0_059_net_fail R0_059_dim_fail R1_059_net_fail R1_059_dim_fail
+ R0_060 R1_060 R0_060_net_fail R0_060_dim_fail R1_060_net_fail R1_060_dim_fail
+ R0_061 R1_061 R0_061_net_fail R0_061_dim_fail R1_061_net_fail R1_061_dim_fail
+ R0_062 R1_062 R0_062_net_fail R0_062_dim_fail R1_062_net_fail R1_062_dim_fail
+ R0_063 R1_063 R0_063_net_fail R0_063_dim_fail R1_063_net_fail R1_063_dim_fail

R000 R0_000 R1_000 sky130_fd_pr__res_xhigh_po_2p85 l=3.35 w=2.85

R001 R0_001 R1_001 sky130_fd_pr__res_xhigh_po_2p85 l=6.7 w=2.85

R002 R0_002 R1_002 sky130_fd_pr__res_xhigh_po_2p85 l=10.05 w=2.85

R003 R0_003 R1_003 sky130_fd_pr__res_xhigh_po_2p85 l=13.4 w=2.85

R004 R0_004 R1_004 sky130_fd_pr__res_xhigh_po_2p85 l=16.75 w=2.85

R005 R0_005 R1_005 sky130_fd_pr__res_xhigh_po_2p85 l=20.1 w=2.85

R006 R0_006 R1_006 sky130_fd_pr__res_xhigh_po_2p85 l=23.45 w=2.85

R007 R0_007 R1_007 sky130_fd_pr__res_xhigh_po_2p85 l=26.8 w=2.85

R008 R0_008 R1_008 sky130_fd_pr__res_xhigh_po_2p85 l=6.7 w=2.85

R009 R0_009 R1_009 sky130_fd_pr__res_xhigh_po_2p85 l=13.4 w=2.85

R010 R0_010 R1_010 sky130_fd_pr__res_xhigh_po_2p85 l=20.1 w=2.85

R011 R0_011 R1_011 sky130_fd_pr__res_xhigh_po_2p85 l=26.8 w=2.85

R012 R0_012 R1_012 sky130_fd_pr__res_xhigh_po_2p85 l=33.5 w=2.85

R013 R0_013 R1_013 sky130_fd_pr__res_xhigh_po_2p85 l=40.2 w=2.85

R014 R0_014 R1_014 sky130_fd_pr__res_xhigh_po_2p85 l=46.9 w=2.85

R015 R0_015 R1_015 sky130_fd_pr__res_xhigh_po_2p85 l=53.6 w=2.85

R016 R0_016 R1_016 sky130_fd_pr__res_xhigh_po_2p85 l=10.05 w=2.85

R017 R0_017 R1_017 sky130_fd_pr__res_xhigh_po_2p85 l=20.1 w=2.85

R018 R0_018 R1_018 sky130_fd_pr__res_xhigh_po_2p85 l=30.15 w=2.85

R019 R0_019 R1_019 sky130_fd_pr__res_xhigh_po_2p85 l=40.2 w=2.85

R020 R0_020 R1_020 sky130_fd_pr__res_xhigh_po_2p85 l=50.25 w=2.85

R021 R0_021 R1_021 sky130_fd_pr__res_xhigh_po_2p85 l=60.3 w=2.85

R022 R0_022 R1_022 sky130_fd_pr__res_xhigh_po_2p85 l=70.35 w=2.85

R023 R0_023 R1_023 sky130_fd_pr__res_xhigh_po_2p85 l=80.4 w=2.85

R024 R0_024 R1_024 sky130_fd_pr__res_xhigh_po_2p85 l=13.4 w=2.85

R025 R0_025 R1_025 sky130_fd_pr__res_xhigh_po_2p85 l=26.8 w=2.85

R026 R0_026 R1_026 sky130_fd_pr__res_xhigh_po_2p85 l=40.2 w=2.85

R027 R0_027 R1_027 sky130_fd_pr__res_xhigh_po_2p85 l=53.6 w=2.85

R028 R0_028 R1_028 sky130_fd_pr__res_xhigh_po_2p85 l=67.0 w=2.85

R029 R0_029 R1_029 sky130_fd_pr__res_xhigh_po_2p85 l=80.4 w=2.85

R030 R0_030 R1_030 sky130_fd_pr__res_xhigh_po_2p85 l=93.8 w=2.85

R031 R0_031 R1_031 sky130_fd_pr__res_xhigh_po_2p85 l=107.2 w=2.85

R032 R0_032 R1_032 sky130_fd_pr__res_xhigh_po_2p85 l=16.75 w=2.85

R033 R0_033 R1_033 sky130_fd_pr__res_xhigh_po_2p85 l=33.5 w=2.85

R034 R0_034 R1_034 sky130_fd_pr__res_xhigh_po_2p85 l=50.25 w=2.85

R035 R0_035 R1_035 sky130_fd_pr__res_xhigh_po_2p85 l=67.0 w=2.85

R036 R0_036 R1_036 sky130_fd_pr__res_xhigh_po_2p85 l=83.75 w=2.85

R037 R0_037 R1_037 sky130_fd_pr__res_xhigh_po_2p85 l=100.5 w=2.85

R038 R0_038 R1_038 sky130_fd_pr__res_xhigh_po_2p85 l=117.25 w=2.85

R039 R0_039 R1_039 sky130_fd_pr__res_xhigh_po_2p85 l=134.0 w=2.85

R040 R0_040 R1_040 sky130_fd_pr__res_xhigh_po_2p85 l=20.1 w=2.85

R041 R0_041 R1_041 sky130_fd_pr__res_xhigh_po_2p85 l=40.2 w=2.85

R042 R0_042 R1_042 sky130_fd_pr__res_xhigh_po_2p85 l=60.3 w=2.85

R043 R0_043 R1_043 sky130_fd_pr__res_xhigh_po_2p85 l=80.4 w=2.85

R044 R0_044 R1_044 sky130_fd_pr__res_xhigh_po_2p85 l=100.5 w=2.85

R045 R0_045 R1_045 sky130_fd_pr__res_xhigh_po_2p85 l=120.6 w=2.85

R046 R0_046 R1_046 sky130_fd_pr__res_xhigh_po_2p85 l=140.7 w=2.85

R047 R0_047 R1_047 sky130_fd_pr__res_xhigh_po_2p85 l=160.8 w=2.85

R048 R0_048 R1_048 sky130_fd_pr__res_xhigh_po_2p85 l=23.45 w=2.85

R049 R0_049 R1_049 sky130_fd_pr__res_xhigh_po_2p85 l=46.9 w=2.85

R050 R0_050 R1_050 sky130_fd_pr__res_xhigh_po_2p85 l=70.35 w=2.85

R051 R0_051 R1_051 sky130_fd_pr__res_xhigh_po_2p85 l=93.8 w=2.85

R052 R0_052 R1_052 sky130_fd_pr__res_xhigh_po_2p85 l=117.25 w=2.85

R053 R0_053 R1_053 sky130_fd_pr__res_xhigh_po_2p85 l=140.7 w=2.85

R054 R0_054 R1_054 sky130_fd_pr__res_xhigh_po_2p85 l=164.15 w=2.85

R055 R0_055 R1_055 sky130_fd_pr__res_xhigh_po_2p85 l=187.6 w=2.85

R056 R0_056 R1_056 sky130_fd_pr__res_xhigh_po_2p85 l=26.8 w=2.85

R057 R0_057 R1_057 sky130_fd_pr__res_xhigh_po_2p85 l=53.6 w=2.85

R058 R0_058 R1_058 sky130_fd_pr__res_xhigh_po_2p85 l=80.4 w=2.85

R059 R0_059 R1_059 sky130_fd_pr__res_xhigh_po_2p85 l=107.2 w=2.85

R060 R0_060 R1_060 sky130_fd_pr__res_xhigh_po_2p85 l=134.0 w=2.85

R061 R0_061 R1_061 sky130_fd_pr__res_xhigh_po_2p85 l=160.8 w=2.85

R062 R0_062 R1_062 sky130_fd_pr__res_xhigh_po_2p85 l=187.6 w=2.85

R063 R0_063 R1_063 sky130_fd_pr__res_xhigh_po_2p85 l=214.4 w=2.85

R000_net_fail R0_000_net_fail R1_000_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=5.025 w=4.275

R001_net_fail R0_001_net_fail R1_001_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=10.05 w=4.275

R002_net_fail R0_002_net_fail R1_002_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=15.075000000000001 w=4.275

R003_net_fail R0_003_net_fail R1_003_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=20.1 w=4.275

R004_net_fail R0_004_net_fail R1_004_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=25.125 w=4.275

R005_net_fail R0_005_net_fail R1_005_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=30.150000000000002 w=4.275

R006_net_fail R0_006_net_fail R1_006_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=35.175 w=4.275

R007_net_fail R0_007_net_fail R1_007_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=40.2 w=4.275

R008_net_fail R0_008_net_fail R1_008_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=10.05 w=4.275

R009_net_fail R0_009_net_fail R1_009_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=20.1 w=4.275

R010_net_fail R0_010_net_fail R1_010_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=30.150000000000002 w=4.275

R011_net_fail R0_011_net_fail R1_011_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=40.2 w=4.275

R012_net_fail R0_012_net_fail R1_012_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=50.25 w=4.275

R013_net_fail R0_013_net_fail R1_013_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=60.300000000000004 w=4.275

R014_net_fail R0_014_net_fail R1_014_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=70.35 w=4.275

R015_net_fail R0_015_net_fail R1_015_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=80.4 w=4.275

R016_net_fail R0_016_net_fail R1_016_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=15.075000000000001 w=4.275

R017_net_fail R0_017_net_fail R1_017_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=30.150000000000002 w=4.275

R018_net_fail R0_018_net_fail R1_018_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=45.224999999999994 w=4.275

R019_net_fail R0_019_net_fail R1_019_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=60.300000000000004 w=4.275

R020_net_fail R0_020_net_fail R1_020_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=75.375 w=4.275

R021_net_fail R0_021_net_fail R1_021_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=90.44999999999999 w=4.275

R022_net_fail R0_022_net_fail R1_022_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=105.52499999999999 w=4.275

R023_net_fail R0_023_net_fail R1_023_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=120.60000000000001 w=4.275

R024_net_fail R0_024_net_fail R1_024_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=20.1 w=4.275

R025_net_fail R0_025_net_fail R1_025_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=40.2 w=4.275

R026_net_fail R0_026_net_fail R1_026_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=60.300000000000004 w=4.275

R027_net_fail R0_027_net_fail R1_027_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=80.4 w=4.275

R028_net_fail R0_028_net_fail R1_028_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=100.5 w=4.275

R029_net_fail R0_029_net_fail R1_029_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=120.60000000000001 w=4.275

R030_net_fail R0_030_net_fail R1_030_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=140.7 w=4.275

R031_net_fail R0_031_net_fail R1_031_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=160.8 w=4.275

R032_net_fail R0_032_net_fail R1_032_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=25.125 w=4.275

R033_net_fail R0_033_net_fail R1_033_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=50.25 w=4.275

R034_net_fail R0_034_net_fail R1_034_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=75.375 w=4.275

R035_net_fail R0_035_net_fail R1_035_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=100.5 w=4.275

R036_net_fail R0_036_net_fail R1_036_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=125.625 w=4.275

R037_net_fail R0_037_net_fail R1_037_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=150.75 w=4.275

R038_net_fail R0_038_net_fail R1_038_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=175.875 w=4.275

R039_net_fail R0_039_net_fail R1_039_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=201.0 w=4.275

R040_net_fail R0_040_net_fail R1_040_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=30.150000000000002 w=4.275

R041_net_fail R0_041_net_fail R1_041_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=60.300000000000004 w=4.275

R042_net_fail R0_042_net_fail R1_042_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=90.44999999999999 w=4.275

R043_net_fail R0_043_net_fail R1_043_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=120.60000000000001 w=4.275

R044_net_fail R0_044_net_fail R1_044_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=150.75 w=4.275

R045_net_fail R0_045_net_fail R1_045_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=180.89999999999998 w=4.275

R046_net_fail R0_046_net_fail R1_046_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=211.04999999999998 w=4.275

R047_net_fail R0_047_net_fail R1_047_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=241.20000000000002 w=4.275

R048_net_fail R0_048_net_fail R1_048_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=35.175 w=4.275

R049_net_fail R0_049_net_fail R1_049_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=70.35 w=4.275

R050_net_fail R0_050_net_fail R1_050_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=105.52499999999999 w=4.275

R051_net_fail R0_051_net_fail R1_051_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=140.7 w=4.275

R052_net_fail R0_052_net_fail R1_052_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=175.875 w=4.275

R053_net_fail R0_053_net_fail R1_053_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=211.04999999999998 w=4.275

R054_net_fail R0_054_net_fail R1_054_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=246.22500000000002 w=4.275

R055_net_fail R0_055_net_fail R1_055_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=281.4 w=4.275

R056_net_fail R0_056_net_fail R1_056_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=40.2 w=4.275

R057_net_fail R0_057_net_fail R1_057_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=80.4 w=4.275

R058_net_fail R0_058_net_fail R1_058_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=120.60000000000001 w=4.275

R059_net_fail R0_059_net_fail R1_059_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=160.8 w=4.275

R060_net_fail R0_060_net_fail R1_060_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=201.0 w=4.275

R061_net_fail R0_061_net_fail R1_061_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=241.20000000000002 w=4.275

R062_net_fail R0_062_net_fail R1_062_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=281.4 w=4.275

R063_net_fail R0_063_net_fail R1_063_net_fail sky130_fd_pr__res_xhigh_po_2p85 l=321.6 w=4.275

R000_dim_fail R0_000_dim_fail R1_000_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=3.35 w=2.85

R001_dim_fail R0_001_dim_fail R1_001_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=6.7 w=2.85

R002_dim_fail R0_002_dim_fail R1_002_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=10.05 w=2.85

R003_dim_fail R0_003_dim_fail R1_003_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=13.4 w=2.85

R004_dim_fail R0_004_dim_fail R1_004_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=16.75 w=2.85

R005_dim_fail R0_005_dim_fail R1_005_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=20.1 w=2.85

R006_dim_fail R0_006_dim_fail R1_006_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=23.45 w=2.85

R007_dim_fail R0_007_dim_fail R1_007_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=26.8 w=2.85

R008_dim_fail R0_008_dim_fail R1_008_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=6.7 w=2.85

R009_dim_fail R0_009_dim_fail R1_009_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=13.4 w=2.85

R010_dim_fail R0_010_dim_fail R1_010_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=20.1 w=2.85

R011_dim_fail R0_011_dim_fail R1_011_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=26.8 w=2.85

R012_dim_fail R0_012_dim_fail R1_012_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=33.5 w=2.85

R013_dim_fail R0_013_dim_fail R1_013_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=40.2 w=2.85

R014_dim_fail R0_014_dim_fail R1_014_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=46.9 w=2.85

R015_dim_fail R0_015_dim_fail R1_015_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=53.6 w=2.85

R016_dim_fail R0_016_dim_fail R1_016_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=10.05 w=2.85

R017_dim_fail R0_017_dim_fail R1_017_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=20.1 w=2.85

R018_dim_fail R0_018_dim_fail R1_018_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=30.15 w=2.85

R019_dim_fail R0_019_dim_fail R1_019_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=40.2 w=2.85

R020_dim_fail R0_020_dim_fail R1_020_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=50.25 w=2.85

R021_dim_fail R0_021_dim_fail R1_021_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=60.3 w=2.85

R022_dim_fail R0_022_dim_fail R1_022_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=70.35 w=2.85

R023_dim_fail R0_023_dim_fail R1_023_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=80.4 w=2.85

R024_dim_fail R0_024_dim_fail R1_024_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=13.4 w=2.85

R025_dim_fail R0_025_dim_fail R1_025_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=26.8 w=2.85

R026_dim_fail R0_026_dim_fail R1_026_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=40.2 w=2.85

R027_dim_fail R0_027_dim_fail R1_027_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=53.6 w=2.85

R028_dim_fail R0_028_dim_fail R1_028_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=67.0 w=2.85

R029_dim_fail R0_029_dim_fail R1_029_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=80.4 w=2.85

R030_dim_fail R0_030_dim_fail R1_030_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=93.8 w=2.85

R031_dim_fail R0_031_dim_fail R1_031_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=107.2 w=2.85

R032_dim_fail R0_032_dim_fail R1_032_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=16.75 w=2.85

R033_dim_fail R0_033_dim_fail R1_033_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=33.5 w=2.85

R034_dim_fail R0_034_dim_fail R1_034_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=50.25 w=2.85

R035_dim_fail R0_035_dim_fail R1_035_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=67.0 w=2.85

R036_dim_fail R0_036_dim_fail R1_036_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=83.75 w=2.85

R037_dim_fail R0_037_dim_fail R1_037_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=100.5 w=2.85

R038_dim_fail R0_038_dim_fail R1_038_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=117.25 w=2.85

R039_dim_fail R0_039_dim_fail R1_039_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=134.0 w=2.85

R040_dim_fail R0_040_dim_fail R1_040_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=20.1 w=2.85

R041_dim_fail R0_041_dim_fail R1_041_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=40.2 w=2.85

R042_dim_fail R0_042_dim_fail R1_042_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=60.3 w=2.85

R043_dim_fail R0_043_dim_fail R1_043_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=80.4 w=2.85

R044_dim_fail R0_044_dim_fail R1_044_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=100.5 w=2.85

R045_dim_fail R0_045_dim_fail R1_045_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=120.6 w=2.85

R046_dim_fail R0_046_dim_fail R1_046_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=140.7 w=2.85

R047_dim_fail R0_047_dim_fail R1_047_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=160.8 w=2.85

R048_dim_fail R0_048_dim_fail R1_048_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=23.45 w=2.85

R049_dim_fail R0_049_dim_fail R1_049_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=46.9 w=2.85

R050_dim_fail R0_050_dim_fail R1_050_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=70.35 w=2.85

R051_dim_fail R0_051_dim_fail R1_051_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=93.8 w=2.85

R052_dim_fail R0_052_dim_fail R1_052_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=117.25 w=2.85

R053_dim_fail R0_053_dim_fail R1_053_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=140.7 w=2.85

R054_dim_fail R0_054_dim_fail R1_054_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=164.15 w=2.85

R055_dim_fail R0_055_dim_fail R1_055_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=187.6 w=2.85

R056_dim_fail R0_056_dim_fail R1_056_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=26.8 w=2.85

R057_dim_fail R0_057_dim_fail R1_057_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=53.6 w=2.85

R058_dim_fail R0_058_dim_fail R1_058_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=80.4 w=2.85

R059_dim_fail R0_059_dim_fail R1_059_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=107.2 w=2.85

R060_dim_fail R0_060_dim_fail R1_060_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=134.0 w=2.85

R061_dim_fail R0_061_dim_fail R1_061_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=160.8 w=2.85

R062_dim_fail R0_062_dim_fail R1_062_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=187.6 w=2.85

R063_dim_fail R0_063_dim_fail R1_063_dim_fail sky130_fd_pr__res_xhigh_po_2p85 l=214.4 w=2.85

.ENDS