* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O
MI98 n0 D net076 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI14 net076 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 db sceb n0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD net076 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net062 s0 net052 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net052 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net51 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net43 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net43 M1 net51 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net061 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net069 s0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 sceb SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net069 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net061 net062 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 db RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net089 net062 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net062 RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net089 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net062 s0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net54 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net54 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 M0 RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net069 s0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net069 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 sceb SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75U l=0.5U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0U l=0.5U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_hvl__sdfrtp_1
