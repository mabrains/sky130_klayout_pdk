* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_lp__fa_m A B CIN VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I CIN:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
MMIN2 COUT majb VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN nmajmid VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj21 nmajmid A VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND B nmajmid VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 A VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 B VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR B pmajmid VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj30 pmajmid CIN majb VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 pmajmid A VPWR VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.42U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_lp__fa_m
