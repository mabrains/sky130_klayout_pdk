 
* Copyright 2022 Mabrains
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Affero General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Affero General Public License for more details.
* 
* You should have received a copy of the GNU Affero General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
.SUBCKT sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p35 DRAIN GATE SOURCE BULK_lyr_fail

Mx_lyr_fail DRAIN_lyr_fail GATE_lyr_fail SOURCE_lyr_fail BULK_lyr_fail sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p35 w=20.0u l=0.35u nf=4 m=1 ad=0.725p as=0.725p pd=6.16u ps=6.16u nrd=0.058 nrs=0.058 sa=0 sb=0 sd=0

.ENDS