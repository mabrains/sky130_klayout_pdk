 
* Copyright 2022 Mabrains
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Affero General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Affero General Public License for more details.
* 
* You should have received a copy of the GNU Affero General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.

.SUBCKT sky130_fd_pr__res_high_po_0p69 
+ R0_000_net_fail R1_000_net_fail
+ R0_001_net_fail R1_001_net_fail
+ R0_002_net_fail R1_002_net_fail
+ R0_003_net_fail R1_003_net_fail
+ R0_004_net_fail R1_004_net_fail
+ R0_005_net_fail R1_005_net_fail
+ R0_006_net_fail R1_006_net_fail
+ R0_007_net_fail R1_007_net_fail
+ R0_008_net_fail R1_008_net_fail
+ R0_009_net_fail R1_009_net_fail
+ R0_010_net_fail R1_010_net_fail
+ R0_011_net_fail R1_011_net_fail
+ R0_012_net_fail R1_012_net_fail
+ R0_013_net_fail R1_013_net_fail
+ R0_014_net_fail R1_014_net_fail
+ R0_015_net_fail R1_015_net_fail
+ R0_016_net_fail R1_016_net_fail
+ R0_017_net_fail R1_017_net_fail
+ R0_018_net_fail R1_018_net_fail
+ R0_019_net_fail R1_019_net_fail
+ R0_020_net_fail R1_020_net_fail
+ R0_021_net_fail R1_021_net_fail
+ R0_022_net_fail R1_022_net_fail
+ R0_023_net_fail R1_023_net_fail
+ R0_024_net_fail R1_024_net_fail
+ R0_025_net_fail R1_025_net_fail
+ R0_026_net_fail R1_026_net_fail
+ R0_027_net_fail R1_027_net_fail
+ R0_028_net_fail R1_028_net_fail
+ R0_029_net_fail R1_029_net_fail
+ R0_030_net_fail R1_030_net_fail
+ R0_031_net_fail R1_031_net_fail
+ R0_032_net_fail R1_032_net_fail
+ R0_033_net_fail R1_033_net_fail
+ R0_034_net_fail R1_034_net_fail
+ R0_035_net_fail R1_035_net_fail
+ R0_036_net_fail R1_036_net_fail
+ R0_037_net_fail R1_037_net_fail
+ R0_038_net_fail R1_038_net_fail
+ R0_039_net_fail R1_039_net_fail
+ R0_040_net_fail R1_040_net_fail
+ R0_041_net_fail R1_041_net_fail
+ R0_042_net_fail R1_042_net_fail
+ R0_043_net_fail R1_043_net_fail
+ R0_044_net_fail R1_044_net_fail
+ R0_045_net_fail R1_045_net_fail
+ R0_046_net_fail R1_046_net_fail
+ R0_047_net_fail R1_047_net_fail
+ R0_048_net_fail R1_048_net_fail
+ R0_049_net_fail R1_049_net_fail
+ R0_050_net_fail R1_050_net_fail
+ R0_051_net_fail R1_051_net_fail
+ R0_052_net_fail R1_052_net_fail
+ R0_053_net_fail R1_053_net_fail
+ R0_054_net_fail R1_054_net_fail
+ R0_055_net_fail R1_055_net_fail
+ R0_056_net_fail R1_056_net_fail
+ R0_057_net_fail R1_057_net_fail
+ R0_058_net_fail R1_058_net_fail
+ R0_059_net_fail R1_059_net_fail
+ R0_060_net_fail R1_060_net_fail
+ R0_061_net_fail R1_061_net_fail
+ R0_062_net_fail R1_062_net_fail
+ R0_063_net_fail R1_063_net_fail

R000_net_fail R0_000_net_fail R1_000_net_fail sky130_fd_pr__res_high_po_0p69 l=1.4690549999999998u w=0.8518049999999999u

R001_net_fail R0_001_net_fail R1_001_net_fail sky130_fd_pr__res_high_po_0p69 l=2.9381099999999996u w=0.8518049999999999u

R002_net_fail R0_002_net_fail R1_002_net_fail sky130_fd_pr__res_high_po_0p69 l=4.407165u w=0.8518049999999999u

R003_net_fail R0_003_net_fail R1_003_net_fail sky130_fd_pr__res_high_po_0p69 l=5.876219999999999u w=0.8518049999999999u

R004_net_fail R0_004_net_fail R1_004_net_fail sky130_fd_pr__res_high_po_0p69 l=7.345275u w=0.8518049999999999u

R005_net_fail R0_005_net_fail R1_005_net_fail sky130_fd_pr__res_high_po_0p69 l=8.81433u w=0.8518049999999999u

R006_net_fail R0_006_net_fail R1_006_net_fail sky130_fd_pr__res_high_po_0p69 l=10.283384999999999u w=0.8518049999999999u

R007_net_fail R0_007_net_fail R1_007_net_fail sky130_fd_pr__res_high_po_0p69 l=11.752439999999998u w=0.8518049999999999u

R008_net_fail R0_008_net_fail R1_008_net_fail sky130_fd_pr__res_high_po_0p69 l=2.9381099999999996u w=0.8518049999999999u

R009_net_fail R0_009_net_fail R1_009_net_fail sky130_fd_pr__res_high_po_0p69 l=5.876219999999999u w=0.8518049999999999u

R010_net_fail R0_010_net_fail R1_010_net_fail sky130_fd_pr__res_high_po_0p69 l=8.81433u w=0.8518049999999999u

R011_net_fail R0_011_net_fail R1_011_net_fail sky130_fd_pr__res_high_po_0p69 l=11.752439999999998u w=0.8518049999999999u

R012_net_fail R0_012_net_fail R1_012_net_fail sky130_fd_pr__res_high_po_0p69 l=14.69055u w=0.8518049999999999u

R013_net_fail R0_013_net_fail R1_013_net_fail sky130_fd_pr__res_high_po_0p69 l=17.62866u w=0.8518049999999999u

R014_net_fail R0_014_net_fail R1_014_net_fail sky130_fd_pr__res_high_po_0p69 l=20.566769999999998u w=0.8518049999999999u

R015_net_fail R0_015_net_fail R1_015_net_fail sky130_fd_pr__res_high_po_0p69 l=23.504879999999996u w=0.8518049999999999u

R016_net_fail R0_016_net_fail R1_016_net_fail sky130_fd_pr__res_high_po_0p69 l=4.407165u w=0.8518049999999999u

R017_net_fail R0_017_net_fail R1_017_net_fail sky130_fd_pr__res_high_po_0p69 l=8.81433u w=0.8518049999999999u

R018_net_fail R0_018_net_fail R1_018_net_fail sky130_fd_pr__res_high_po_0p69 l=13.221495u w=0.8518049999999999u

R019_net_fail R0_019_net_fail R1_019_net_fail sky130_fd_pr__res_high_po_0p69 l=17.62866u w=0.8518049999999999u

R020_net_fail R0_020_net_fail R1_020_net_fail sky130_fd_pr__res_high_po_0p69 l=22.035825u w=0.8518049999999999u

R021_net_fail R0_021_net_fail R1_021_net_fail sky130_fd_pr__res_high_po_0p69 l=26.44299u w=0.8518049999999999u

R022_net_fail R0_022_net_fail R1_022_net_fail sky130_fd_pr__res_high_po_0p69 l=30.850154999999997u w=0.8518049999999999u

R023_net_fail R0_023_net_fail R1_023_net_fail sky130_fd_pr__res_high_po_0p69 l=35.25732u w=0.8518049999999999u

R024_net_fail R0_024_net_fail R1_024_net_fail sky130_fd_pr__res_high_po_0p69 l=5.876219999999999u w=0.8518049999999999u

R025_net_fail R0_025_net_fail R1_025_net_fail sky130_fd_pr__res_high_po_0p69 l=11.752439999999998u w=0.8518049999999999u

R026_net_fail R0_026_net_fail R1_026_net_fail sky130_fd_pr__res_high_po_0p69 l=17.62866u w=0.8518049999999999u

R027_net_fail R0_027_net_fail R1_027_net_fail sky130_fd_pr__res_high_po_0p69 l=23.504879999999996u w=0.8518049999999999u

R028_net_fail R0_028_net_fail R1_028_net_fail sky130_fd_pr__res_high_po_0p69 l=29.3811u w=0.8518049999999999u

R029_net_fail R0_029_net_fail R1_029_net_fail sky130_fd_pr__res_high_po_0p69 l=35.25732u w=0.8518049999999999u

R030_net_fail R0_030_net_fail R1_030_net_fail sky130_fd_pr__res_high_po_0p69 l=41.133539999999996u w=0.8518049999999999u

R031_net_fail R0_031_net_fail R1_031_net_fail sky130_fd_pr__res_high_po_0p69 l=47.00975999999999u w=0.8518049999999999u

R032_net_fail R0_032_net_fail R1_032_net_fail sky130_fd_pr__res_high_po_0p69 l=7.345275u w=0.8518049999999999u

R033_net_fail R0_033_net_fail R1_033_net_fail sky130_fd_pr__res_high_po_0p69 l=14.69055u w=0.8518049999999999u

R034_net_fail R0_034_net_fail R1_034_net_fail sky130_fd_pr__res_high_po_0p69 l=22.035825u w=0.8518049999999999u

R035_net_fail R0_035_net_fail R1_035_net_fail sky130_fd_pr__res_high_po_0p69 l=29.3811u w=0.8518049999999999u

R036_net_fail R0_036_net_fail R1_036_net_fail sky130_fd_pr__res_high_po_0p69 l=36.726375u w=0.8518049999999999u

R037_net_fail R0_037_net_fail R1_037_net_fail sky130_fd_pr__res_high_po_0p69 l=44.07165u w=0.8518049999999999u

R038_net_fail R0_038_net_fail R1_038_net_fail sky130_fd_pr__res_high_po_0p69 l=51.41692499999999u w=0.8518049999999999u

R039_net_fail R0_039_net_fail R1_039_net_fail sky130_fd_pr__res_high_po_0p69 l=58.7622u w=0.8518049999999999u

R040_net_fail R0_040_net_fail R1_040_net_fail sky130_fd_pr__res_high_po_0p69 l=8.81433u w=0.8518049999999999u

R041_net_fail R0_041_net_fail R1_041_net_fail sky130_fd_pr__res_high_po_0p69 l=17.62866u w=0.8518049999999999u

R042_net_fail R0_042_net_fail R1_042_net_fail sky130_fd_pr__res_high_po_0p69 l=26.44299u w=0.8518049999999999u

R043_net_fail R0_043_net_fail R1_043_net_fail sky130_fd_pr__res_high_po_0p69 l=35.25732u w=0.8518049999999999u

R044_net_fail R0_044_net_fail R1_044_net_fail sky130_fd_pr__res_high_po_0p69 l=44.07165u w=0.8518049999999999u

R045_net_fail R0_045_net_fail R1_045_net_fail sky130_fd_pr__res_high_po_0p69 l=52.88598u w=0.8518049999999999u

R046_net_fail R0_046_net_fail R1_046_net_fail sky130_fd_pr__res_high_po_0p69 l=61.700309999999995u w=0.8518049999999999u

R047_net_fail R0_047_net_fail R1_047_net_fail sky130_fd_pr__res_high_po_0p69 l=70.51464u w=0.8518049999999999u

R048_net_fail R0_048_net_fail R1_048_net_fail sky130_fd_pr__res_high_po_0p69 l=10.283384999999999u w=0.8518049999999999u

R049_net_fail R0_049_net_fail R1_049_net_fail sky130_fd_pr__res_high_po_0p69 l=20.566769999999998u w=0.8518049999999999u

R050_net_fail R0_050_net_fail R1_050_net_fail sky130_fd_pr__res_high_po_0p69 l=30.850154999999997u w=0.8518049999999999u

R051_net_fail R0_051_net_fail R1_051_net_fail sky130_fd_pr__res_high_po_0p69 l=41.133539999999996u w=0.8518049999999999u

R052_net_fail R0_052_net_fail R1_052_net_fail sky130_fd_pr__res_high_po_0p69 l=51.41692499999999u w=0.8518049999999999u

R053_net_fail R0_053_net_fail R1_053_net_fail sky130_fd_pr__res_high_po_0p69 l=61.700309999999995u w=0.8518049999999999u

R054_net_fail R0_054_net_fail R1_054_net_fail sky130_fd_pr__res_high_po_0p69 l=71.983695u w=0.8518049999999999u

R055_net_fail R0_055_net_fail R1_055_net_fail sky130_fd_pr__res_high_po_0p69 l=82.26707999999999u w=0.8518049999999999u

R056_net_fail R0_056_net_fail R1_056_net_fail sky130_fd_pr__res_high_po_0p69 l=11.752439999999998u w=0.8518049999999999u

R057_net_fail R0_057_net_fail R1_057_net_fail sky130_fd_pr__res_high_po_0p69 l=23.504879999999996u w=0.8518049999999999u

R058_net_fail R0_058_net_fail R1_058_net_fail sky130_fd_pr__res_high_po_0p69 l=35.25732u w=0.8518049999999999u

R059_net_fail R0_059_net_fail R1_059_net_fail sky130_fd_pr__res_high_po_0p69 l=47.00975999999999u w=0.8518049999999999u

R060_net_fail R0_060_net_fail R1_060_net_fail sky130_fd_pr__res_high_po_0p69 l=58.7622u w=0.8518049999999999u

R061_net_fail R0_061_net_fail R1_061_net_fail sky130_fd_pr__res_high_po_0p69 l=70.51464u w=0.8518049999999999u

R062_net_fail R0_062_net_fail R1_062_net_fail sky130_fd_pr__res_high_po_0p69 l=82.26707999999999u w=0.8518049999999999u

R063_net_fail R0_063_net_fail R1_063_net_fail sky130_fd_pr__res_high_po_0p69 l=94.01951999999999u w=0.8518049999999999u

.ENDS