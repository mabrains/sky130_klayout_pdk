* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.subckt_dim_fail sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1m5_floatm4_top C0_dim_fail C1_dim_fail M5_dim_fail SUB

Csky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1m5_floatm4_0[0|0] M5_dim_fail C1_dim_fail C0_dim_fail SUB sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1m5_floatm4

Csky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1m5_floatm4_0[1|0] M5_dim_fail C1_dim_fail C0_dim_fail SUB sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1m5_floatm4

Csky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1m5_floatm4_0[0|1] M5_dim_fail C1_dim_fail C0_dim_fail SUB sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1m5_floatm4

Csky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1m5_floatm4_0[1|1] M5_dim_fail C1_dim_fail C0_dim_fail SUB sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1m5_floatm4

.ends_dim_fail

.ENDS