 
* Copyright 2022 SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT connectivity_m4 SUB_SRC_D1 GAT_DRN_R0 D0_R1

M0 SUB_SRC_D1 GAT_DRN_R0 GAT_DRN_R0 SUB_SRC_D1 sky130_fd_pr__nfet_01v8 w=0.42U l=0.15U nf=1

D0 D0_R1 SUB_SRC_D1 sky130_fd_pr__diode_pd2nw_05v5 A=0.2025P P=1.8U

R0 GAT_DRN_R0 D0_R1 SUB_SRC_D1 sky130_fd_pr__res_generic_nd l=2.1U w=0.42U

.ENDS
