* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3 C0 C1 SUB MET3
*.PININFO C0:? C1:? SUB:? MET3:?
+ sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3_dim_fail

C1_dim_fail C0_dim_fail C1_dim_fail SUB MET3_dim_fail

.ENDS