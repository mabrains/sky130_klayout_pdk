 
* Copyright 2022 Mabrains
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Affero General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Affero General Public License for more details.
* 
* You should have received a copy of the GNU Affero General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
.SUBCKT sky130_fd_pr__rf_pfet_01v8_aF08W1p68L0p15 DRAIN GATE SOURCE BULK_lyr_fail

Mx_lyr_fail DRAIN_lyr_fail GATE_lyr_fail SOURCE_lyr_fail BULK_lyr_fail sky130_fd_pr__rf_pfet_01v8_aF08W1p68L0p15 w=13.44u l=0.15u nf=8 m=1 ad=0.2436p as=0.2436p pd=4.0u ps=4.0u nrd=0.1726 nrs=0.1726 sa=0 sb=0 sd=0

.ENDS