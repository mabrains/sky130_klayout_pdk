 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__diode_pd2nw_05v5
+ D0_000 D1_000 D0_000_net_fail D0_000_dim_fail D1_000_net_fail D1_000_dim_fail
+ D0_001 D1_001 D0_001_net_fail D0_001_dim_fail D1_001_net_fail D1_001_dim_fail
+ D0_002 D1_002 D0_002_net_fail D0_002_dim_fail D1_002_net_fail D1_002_dim_fail
+ D0_003 D1_003 D0_003_net_fail D0_003_dim_fail D1_003_net_fail D1_003_dim_fail
+ D0_004 D1_004 D0_004_net_fail D0_004_dim_fail D1_004_net_fail D1_004_dim_fail
+ D0_005 D1_005 D0_005_net_fail D0_005_dim_fail D1_005_net_fail D1_005_dim_fail
+ D0_006 D1_006 D0_006_net_fail D0_006_dim_fail D1_006_net_fail D1_006_dim_fail
+ D0_007 D1_007 D0_007_net_fail D0_007_dim_fail D1_007_net_fail D1_007_dim_fail
+ D0_008 D1_008 D0_008_net_fail D0_008_dim_fail D1_008_net_fail D1_008_dim_fail
+ D0_009 D1_009 D0_009_net_fail D0_009_dim_fail D1_009_net_fail D1_009_dim_fail
+ D0_010 D1_010 D0_010_net_fail D0_010_dim_fail D1_010_net_fail D1_010_dim_fail
+ D0_011 D1_011 D0_011_net_fail D0_011_dim_fail D1_011_net_fail D1_011_dim_fail
+ D0_012 D1_012 D0_012_net_fail D0_012_dim_fail D1_012_net_fail D1_012_dim_fail
+ D0_013 D1_013 D0_013_net_fail D0_013_dim_fail D1_013_net_fail D1_013_dim_fail
+ D0_014 D1_014 D0_014_net_fail D0_014_dim_fail D1_014_net_fail D1_014_dim_fail
+ D0_015 D1_015 D0_015_net_fail D0_015_dim_fail D1_015_net_fail D1_015_dim_fail
+ D0_016 D1_016 D0_016_net_fail D0_016_dim_fail D1_016_net_fail D1_016_dim_fail
+ D0_017 D1_017 D0_017_net_fail D0_017_dim_fail D1_017_net_fail D1_017_dim_fail
+ D0_018 D1_018 D0_018_net_fail D0_018_dim_fail D1_018_net_fail D1_018_dim_fail
+ D0_019 D1_019 D0_019_net_fail D0_019_dim_fail D1_019_net_fail D1_019_dim_fail
+ D0_020 D1_020 D0_020_net_fail D0_020_dim_fail D1_020_net_fail D1_020_dim_fail
+ D0_021 D1_021 D0_021_net_fail D0_021_dim_fail D1_021_net_fail D1_021_dim_fail
+ D0_022 D1_022 D0_022_net_fail D0_022_dim_fail D1_022_net_fail D1_022_dim_fail
+ D0_023 D1_023 D0_023_net_fail D0_023_dim_fail D1_023_net_fail D1_023_dim_fail
+ D0_024 D1_024 D0_024_net_fail D0_024_dim_fail D1_024_net_fail D1_024_dim_fail
+ D0_025 D1_025 D0_025_net_fail D0_025_dim_fail D1_025_net_fail D1_025_dim_fail
+ D0_026 D1_026 D0_026_net_fail D0_026_dim_fail D1_026_net_fail D1_026_dim_fail
+ D0_027 D1_027 D0_027_net_fail D0_027_dim_fail D1_027_net_fail D1_027_dim_fail
+ D0_028 D1_028 D0_028_net_fail D0_028_dim_fail D1_028_net_fail D1_028_dim_fail
+ D0_029 D1_029 D0_029_net_fail D0_029_dim_fail D1_029_net_fail D1_029_dim_fail
+ D0_030 D1_030 D0_030_net_fail D0_030_dim_fail D1_030_net_fail D1_030_dim_fail
+ D0_031 D1_031 D0_031_net_fail D0_031_dim_fail D1_031_net_fail D1_031_dim_fail
+ D0_032 D1_032 D0_032_net_fail D0_032_dim_fail D1_032_net_fail D1_032_dim_fail
+ D0_033 D1_033 D0_033_net_fail D0_033_dim_fail D1_033_net_fail D1_033_dim_fail
+ D0_034 D1_034 D0_034_net_fail D0_034_dim_fail D1_034_net_fail D1_034_dim_fail
+ D0_035 D1_035 D0_035_net_fail D0_035_dim_fail D1_035_net_fail D1_035_dim_fail
+ D0_036 D1_036 D0_036_net_fail D0_036_dim_fail D1_036_net_fail D1_036_dim_fail
+ D0_037 D1_037 D0_037_net_fail D0_037_dim_fail D1_037_net_fail D1_037_dim_fail
+ D0_038 D1_038 D0_038_net_fail D0_038_dim_fail D1_038_net_fail D1_038_dim_fail
+ D0_039 D1_039 D0_039_net_fail D0_039_dim_fail D1_039_net_fail D1_039_dim_fail
+ D0_040 D1_040 D0_040_net_fail D0_040_dim_fail D1_040_net_fail D1_040_dim_fail
+ D0_041 D1_041 D0_041_net_fail D0_041_dim_fail D1_041_net_fail D1_041_dim_fail
+ D0_042 D1_042 D0_042_net_fail D0_042_dim_fail D1_042_net_fail D1_042_dim_fail
+ D0_043 D1_043 D0_043_net_fail D0_043_dim_fail D1_043_net_fail D1_043_dim_fail
+ D0_044 D1_044 D0_044_net_fail D0_044_dim_fail D1_044_net_fail D1_044_dim_fail
+ D0_045 D1_045 D0_045_net_fail D0_045_dim_fail D1_045_net_fail D1_045_dim_fail
+ D0_046 D1_046 D0_046_net_fail D0_046_dim_fail D1_046_net_fail D1_046_dim_fail
+ D0_047 D1_047 D0_047_net_fail D0_047_dim_fail D1_047_net_fail D1_047_dim_fail
+ D0_048 D1_048 D0_048_net_fail D0_048_dim_fail D1_048_net_fail D1_048_dim_fail
+ D0_049 D1_049 D0_049_net_fail D0_049_dim_fail D1_049_net_fail D1_049_dim_fail
+ D0_050 D1_050 D0_050_net_fail D0_050_dim_fail D1_050_net_fail D1_050_dim_fail
+ D0_051 D1_051 D0_051_net_fail D0_051_dim_fail D1_051_net_fail D1_051_dim_fail
+ D0_052 D1_052 D0_052_net_fail D0_052_dim_fail D1_052_net_fail D1_052_dim_fail
+ D0_053 D1_053 D0_053_net_fail D0_053_dim_fail D1_053_net_fail D1_053_dim_fail
+ D0_054 D1_054 D0_054_net_fail D0_054_dim_fail D1_054_net_fail D1_054_dim_fail
+ D0_055 D1_055 D0_055_net_fail D0_055_dim_fail D1_055_net_fail D1_055_dim_fail
+ D0_056 D1_056 D0_056_net_fail D0_056_dim_fail D1_056_net_fail D1_056_dim_fail
+ D0_057 D1_057 D0_057_net_fail D0_057_dim_fail D1_057_net_fail D1_057_dim_fail
+ D0_058 D1_058 D0_058_net_fail D0_058_dim_fail D1_058_net_fail D1_058_dim_fail
+ D0_059 D1_059 D0_059_net_fail D0_059_dim_fail D1_059_net_fail D1_059_dim_fail
+ D0_060 D1_060 D0_060_net_fail D0_060_dim_fail D1_060_net_fail D1_060_dim_fail
+ D0_061 D1_061 D0_061_net_fail D0_061_dim_fail D1_061_net_fail D1_061_dim_fail
+ D0_062 D1_062 D0_062_net_fail D0_062_dim_fail D1_062_net_fail D1_062_dim_fail
+ D0_063 D1_063 D0_063_net_fail D0_063_dim_fail D1_063_net_fail D1_063_dim_fail

D000 D0_000 D1_000 sky130_fd_pr__diode_pd2nw_05v5 AREA=0.2025 PJ=1.8

D001 D0_001 D1_001 sky130_fd_pr__diode_pd2nw_05v5 AREA=0.405 PJ=2.7

D002 D0_002 D1_002 sky130_fd_pr__diode_pd2nw_05v5 AREA=0.6075 PJ=3.6

D003 D0_003 D1_003 sky130_fd_pr__diode_pd2nw_05v5 AREA=0.81 PJ=4.5

D004 D0_004 D1_004 sky130_fd_pr__diode_pd2nw_05v5 AREA=1.0125 PJ=5.4

D005 D0_005 D1_005 sky130_fd_pr__diode_pd2nw_05v5 AREA=1.215 PJ=6.3

D006 D0_006 D1_006 sky130_fd_pr__diode_pd2nw_05v5 AREA=1.4175 PJ=7.2

D007 D0_007 D1_007 sky130_fd_pr__diode_pd2nw_05v5 AREA=1.62 PJ=8.1

D008 D0_008 D1_008 sky130_fd_pr__diode_pd2nw_05v5 AREA=0.405 PJ=2.7

D009 D0_009 D1_009 sky130_fd_pr__diode_pd2nw_05v5 AREA=0.81 PJ=3.6

D010 D0_010 D1_010 sky130_fd_pr__diode_pd2nw_05v5 AREA=1.215 PJ=4.5

D011 D0_011 D1_011 sky130_fd_pr__diode_pd2nw_05v5 AREA=1.62 PJ=5.4

D012 D0_012 D1_012 sky130_fd_pr__diode_pd2nw_05v5 AREA=2.025 PJ=6.3

D013 D0_013 D1_013 sky130_fd_pr__diode_pd2nw_05v5 AREA=2.43 PJ=7.2

D014 D0_014 D1_014 sky130_fd_pr__diode_pd2nw_05v5 AREA=2.835 PJ=8.1

D015 D0_015 D1_015 sky130_fd_pr__diode_pd2nw_05v5 AREA=3.24 PJ=9.0

D016 D0_016 D1_016 sky130_fd_pr__diode_pd2nw_05v5 AREA=0.6075 PJ=3.6

D017 D0_017 D1_017 sky130_fd_pr__diode_pd2nw_05v5 AREA=1.215 PJ=4.5

D018 D0_018 D1_018 sky130_fd_pr__diode_pd2nw_05v5 AREA=1.8225 PJ=5.4

D019 D0_019 D1_019 sky130_fd_pr__diode_pd2nw_05v5 AREA=2.43 PJ=6.3

D020 D0_020 D1_020 sky130_fd_pr__diode_pd2nw_05v5 AREA=3.0375 PJ=7.2

D021 D0_021 D1_021 sky130_fd_pr__diode_pd2nw_05v5 AREA=3.645 PJ=8.1

D022 D0_022 D1_022 sky130_fd_pr__diode_pd2nw_05v5 AREA=4.2525 PJ=9.0

D023 D0_023 D1_023 sky130_fd_pr__diode_pd2nw_05v5 AREA=4.86 PJ=9.9

D024 D0_024 D1_024 sky130_fd_pr__diode_pd2nw_05v5 AREA=0.81 PJ=4.5

D025 D0_025 D1_025 sky130_fd_pr__diode_pd2nw_05v5 AREA=1.62 PJ=5.4

D026 D0_026 D1_026 sky130_fd_pr__diode_pd2nw_05v5 AREA=2.43 PJ=6.3

D027 D0_027 D1_027 sky130_fd_pr__diode_pd2nw_05v5 AREA=3.24 PJ=7.2

D028 D0_028 D1_028 sky130_fd_pr__diode_pd2nw_05v5 AREA=4.05 PJ=8.1

D029 D0_029 D1_029 sky130_fd_pr__diode_pd2nw_05v5 AREA=4.86 PJ=9.0

D030 D0_030 D1_030 sky130_fd_pr__diode_pd2nw_05v5 AREA=5.67 PJ=9.9

D031 D0_031 D1_031 sky130_fd_pr__diode_pd2nw_05v5 AREA=6.48 PJ=10.8

D032 D0_032 D1_032 sky130_fd_pr__diode_pd2nw_05v5 AREA=1.0125 PJ=5.4

D033 D0_033 D1_033 sky130_fd_pr__diode_pd2nw_05v5 AREA=2.025 PJ=6.3

D034 D0_034 D1_034 sky130_fd_pr__diode_pd2nw_05v5 AREA=3.0375 PJ=7.2

D035 D0_035 D1_035 sky130_fd_pr__diode_pd2nw_05v5 AREA=4.05 PJ=8.1

D036 D0_036 D1_036 sky130_fd_pr__diode_pd2nw_05v5 AREA=5.0625 PJ=9.0

D037 D0_037 D1_037 sky130_fd_pr__diode_pd2nw_05v5 AREA=6.075 PJ=9.9

D038 D0_038 D1_038 sky130_fd_pr__diode_pd2nw_05v5 AREA=7.0875 PJ=10.8

D039 D0_039 D1_039 sky130_fd_pr__diode_pd2nw_05v5 AREA=8.1 PJ=11.7

D040 D0_040 D1_040 sky130_fd_pr__diode_pd2nw_05v5 AREA=1.215 PJ=6.3

D041 D0_041 D1_041 sky130_fd_pr__diode_pd2nw_05v5 AREA=2.43 PJ=7.2

D042 D0_042 D1_042 sky130_fd_pr__diode_pd2nw_05v5 AREA=3.645 PJ=8.1

D043 D0_043 D1_043 sky130_fd_pr__diode_pd2nw_05v5 AREA=4.86 PJ=9.0

D044 D0_044 D1_044 sky130_fd_pr__diode_pd2nw_05v5 AREA=6.075 PJ=9.9

D045 D0_045 D1_045 sky130_fd_pr__diode_pd2nw_05v5 AREA=7.29 PJ=10.8

D046 D0_046 D1_046 sky130_fd_pr__diode_pd2nw_05v5 AREA=8.505 PJ=11.7

D047 D0_047 D1_047 sky130_fd_pr__diode_pd2nw_05v5 AREA=9.72 PJ=12.6

D048 D0_048 D1_048 sky130_fd_pr__diode_pd2nw_05v5 AREA=1.4175 PJ=7.2

D049 D0_049 D1_049 sky130_fd_pr__diode_pd2nw_05v5 AREA=2.835 PJ=8.1

D050 D0_050 D1_050 sky130_fd_pr__diode_pd2nw_05v5 AREA=4.2525 PJ=9.0

D051 D0_051 D1_051 sky130_fd_pr__diode_pd2nw_05v5 AREA=5.67 PJ=9.9

D052 D0_052 D1_052 sky130_fd_pr__diode_pd2nw_05v5 AREA=7.0875 PJ=10.8

D053 D0_053 D1_053 sky130_fd_pr__diode_pd2nw_05v5 AREA=8.505 PJ=11.7

D054 D0_054 D1_054 sky130_fd_pr__diode_pd2nw_05v5 AREA=9.9225 PJ=12.6

D055 D0_055 D1_055 sky130_fd_pr__diode_pd2nw_05v5 AREA=11.34 PJ=13.5

D056 D0_056 D1_056 sky130_fd_pr__diode_pd2nw_05v5 AREA=1.62 PJ=8.1

D057 D0_057 D1_057 sky130_fd_pr__diode_pd2nw_05v5 AREA=3.24 PJ=9.0

D058 D0_058 D1_058 sky130_fd_pr__diode_pd2nw_05v5 AREA=4.86 PJ=9.9

D059 D0_059 D1_059 sky130_fd_pr__diode_pd2nw_05v5 AREA=6.48 PJ=10.8

D060 D0_060 D1_060 sky130_fd_pr__diode_pd2nw_05v5 AREA=8.1 PJ=11.7

D061 D0_061 D1_061 sky130_fd_pr__diode_pd2nw_05v5 AREA=9.72 PJ=12.6

D062 D0_062 D1_062 sky130_fd_pr__diode_pd2nw_05v5 AREA=11.34 PJ=13.5

D063 D0_063 D1_063 sky130_fd_pr__diode_pd2nw_05v5 AREA=12.96 PJ=14.4

D000_net_fail D0_000_net_fail D1_000_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=0.30375 PJ=2.7

D001_net_fail D0_001_net_fail D1_001_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=0.6075 PJ=4.050000000000001

D002_net_fail D0_002_net_fail D1_002_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=0.9112500000000001 PJ=5.4

D003_net_fail D0_003_net_fail D1_003_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.215 PJ=6.75

D004_net_fail D0_004_net_fail D1_004_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.5187499999999998 PJ=8.100000000000001

D005_net_fail D0_005_net_fail D1_005_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.8225000000000002 PJ=9.45

D006_net_fail D0_006_net_fail D1_006_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=2.1262499999999998 PJ=10.8

D007_net_fail D0_007_net_fail D1_007_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=2.43 PJ=12.149999999999999

D008_net_fail D0_008_net_fail D1_008_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=0.6075 PJ=4.050000000000001

D009_net_fail D0_009_net_fail D1_009_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.215 PJ=5.4

D010_net_fail D0_010_net_fail D1_010_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.8225000000000002 PJ=6.75

D011_net_fail D0_011_net_fail D1_011_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=2.43 PJ=8.100000000000001

D012_net_fail D0_012_net_fail D1_012_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=3.0374999999999996 PJ=9.45

D013_net_fail D0_013_net_fail D1_013_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=3.6450000000000005 PJ=10.8

D014_net_fail D0_014_net_fail D1_014_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=4.2524999999999995 PJ=12.149999999999999

D015_net_fail D0_015_net_fail D1_015_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=4.86 PJ=13.5

D016_net_fail D0_016_net_fail D1_016_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=0.9112500000000001 PJ=5.4

D017_net_fail D0_017_net_fail D1_017_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.8225000000000002 PJ=6.75

D018_net_fail D0_018_net_fail D1_018_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=2.73375 PJ=8.100000000000001

D019_net_fail D0_019_net_fail D1_019_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=3.6450000000000005 PJ=9.45

D020_net_fail D0_020_net_fail D1_020_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=4.55625 PJ=10.8

D021_net_fail D0_021_net_fail D1_021_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=5.4675 PJ=12.149999999999999

D022_net_fail D0_022_net_fail D1_022_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=6.37875 PJ=13.5

D023_net_fail D0_023_net_fail D1_023_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=7.290000000000001 PJ=14.850000000000001

D024_net_fail D0_024_net_fail D1_024_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.215 PJ=6.75

D025_net_fail D0_025_net_fail D1_025_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=2.43 PJ=8.100000000000001

D026_net_fail D0_026_net_fail D1_026_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=3.6450000000000005 PJ=9.45

D027_net_fail D0_027_net_fail D1_027_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=4.86 PJ=10.8

D028_net_fail D0_028_net_fail D1_028_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=6.074999999999999 PJ=12.149999999999999

D029_net_fail D0_029_net_fail D1_029_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=7.290000000000001 PJ=13.5

D030_net_fail D0_030_net_fail D1_030_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=8.504999999999999 PJ=14.850000000000001

D031_net_fail D0_031_net_fail D1_031_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=9.72 PJ=16.200000000000003

D032_net_fail D0_032_net_fail D1_032_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.5187499999999998 PJ=8.100000000000001

D033_net_fail D0_033_net_fail D1_033_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=3.0374999999999996 PJ=9.45

D034_net_fail D0_034_net_fail D1_034_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=4.55625 PJ=10.8

D035_net_fail D0_035_net_fail D1_035_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=6.074999999999999 PJ=12.149999999999999

D036_net_fail D0_036_net_fail D1_036_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=7.59375 PJ=13.5

D037_net_fail D0_037_net_fail D1_037_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=9.1125 PJ=14.850000000000001

D038_net_fail D0_038_net_fail D1_038_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=10.631250000000001 PJ=16.200000000000003

D039_net_fail D0_039_net_fail D1_039_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=12.149999999999999 PJ=17.549999999999997

D040_net_fail D0_040_net_fail D1_040_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.8225000000000002 PJ=9.45

D041_net_fail D0_041_net_fail D1_041_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=3.6450000000000005 PJ=10.8

D042_net_fail D0_042_net_fail D1_042_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=5.4675 PJ=12.149999999999999

D043_net_fail D0_043_net_fail D1_043_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=7.290000000000001 PJ=13.5

D044_net_fail D0_044_net_fail D1_044_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=9.1125 PJ=14.850000000000001

D045_net_fail D0_045_net_fail D1_045_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=10.935 PJ=16.200000000000003

D046_net_fail D0_046_net_fail D1_046_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=12.7575 PJ=17.549999999999997

D047_net_fail D0_047_net_fail D1_047_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=14.580000000000002 PJ=18.9

D048_net_fail D0_048_net_fail D1_048_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=2.1262499999999998 PJ=10.8

D049_net_fail D0_049_net_fail D1_049_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=4.2524999999999995 PJ=12.149999999999999

D050_net_fail D0_050_net_fail D1_050_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=6.37875 PJ=13.5

D051_net_fail D0_051_net_fail D1_051_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=8.504999999999999 PJ=14.850000000000001

D052_net_fail D0_052_net_fail D1_052_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=10.631250000000001 PJ=16.200000000000003

D053_net_fail D0_053_net_fail D1_053_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=12.7575 PJ=17.549999999999997

D054_net_fail D0_054_net_fail D1_054_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=14.88375 PJ=18.9

D055_net_fail D0_055_net_fail D1_055_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=17.009999999999998 PJ=20.25

D056_net_fail D0_056_net_fail D1_056_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=2.43 PJ=12.149999999999999

D057_net_fail D0_057_net_fail D1_057_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=4.86 PJ=13.5

D058_net_fail D0_058_net_fail D1_058_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=7.290000000000001 PJ=14.850000000000001

D059_net_fail D0_059_net_fail D1_059_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=9.72 PJ=16.200000000000003

D060_net_fail D0_060_net_fail D1_060_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=12.149999999999999 PJ=17.549999999999997

D061_net_fail D0_061_net_fail D1_061_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=14.580000000000002 PJ=18.9

D062_net_fail D0_062_net_fail D1_062_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=17.009999999999998 PJ=20.25

D063_net_fail D0_063_net_fail D1_063_net_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=19.44 PJ=21.6

D000_dim_fail D0_000_dim_fail D1_000_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=0.2025 PJ=1.8

D001_dim_fail D0_001_dim_fail D1_001_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=0.405 PJ=2.7

D002_dim_fail D0_002_dim_fail D1_002_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=0.6075 PJ=3.6

D003_dim_fail D0_003_dim_fail D1_003_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=0.81 PJ=4.5

D004_dim_fail D0_004_dim_fail D1_004_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.0125 PJ=5.4

D005_dim_fail D0_005_dim_fail D1_005_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.215 PJ=6.3

D006_dim_fail D0_006_dim_fail D1_006_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.4175 PJ=7.2

D007_dim_fail D0_007_dim_fail D1_007_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.62 PJ=8.1

D008_dim_fail D0_008_dim_fail D1_008_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=0.405 PJ=2.7

D009_dim_fail D0_009_dim_fail D1_009_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=0.81 PJ=3.6

D010_dim_fail D0_010_dim_fail D1_010_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.215 PJ=4.5

D011_dim_fail D0_011_dim_fail D1_011_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.62 PJ=5.4

D012_dim_fail D0_012_dim_fail D1_012_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=2.025 PJ=6.3

D013_dim_fail D0_013_dim_fail D1_013_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=2.43 PJ=7.2

D014_dim_fail D0_014_dim_fail D1_014_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=2.835 PJ=8.1

D015_dim_fail D0_015_dim_fail D1_015_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=3.24 PJ=9.0

D016_dim_fail D0_016_dim_fail D1_016_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=0.6075 PJ=3.6

D017_dim_fail D0_017_dim_fail D1_017_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.215 PJ=4.5

D018_dim_fail D0_018_dim_fail D1_018_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.8225 PJ=5.4

D019_dim_fail D0_019_dim_fail D1_019_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=2.43 PJ=6.3

D020_dim_fail D0_020_dim_fail D1_020_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=3.0375 PJ=7.2

D021_dim_fail D0_021_dim_fail D1_021_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=3.645 PJ=8.1

D022_dim_fail D0_022_dim_fail D1_022_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=4.2525 PJ=9.0

D023_dim_fail D0_023_dim_fail D1_023_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=4.86 PJ=9.9

D024_dim_fail D0_024_dim_fail D1_024_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=0.81 PJ=4.5

D025_dim_fail D0_025_dim_fail D1_025_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.62 PJ=5.4

D026_dim_fail D0_026_dim_fail D1_026_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=2.43 PJ=6.3

D027_dim_fail D0_027_dim_fail D1_027_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=3.24 PJ=7.2

D028_dim_fail D0_028_dim_fail D1_028_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=4.05 PJ=8.1

D029_dim_fail D0_029_dim_fail D1_029_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=4.86 PJ=9.0

D030_dim_fail D0_030_dim_fail D1_030_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=5.67 PJ=9.9

D031_dim_fail D0_031_dim_fail D1_031_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=6.48 PJ=10.8

D032_dim_fail D0_032_dim_fail D1_032_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.0125 PJ=5.4

D033_dim_fail D0_033_dim_fail D1_033_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=2.025 PJ=6.3

D034_dim_fail D0_034_dim_fail D1_034_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=3.0375 PJ=7.2

D035_dim_fail D0_035_dim_fail D1_035_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=4.05 PJ=8.1

D036_dim_fail D0_036_dim_fail D1_036_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=5.0625 PJ=9.0

D037_dim_fail D0_037_dim_fail D1_037_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=6.075 PJ=9.9

D038_dim_fail D0_038_dim_fail D1_038_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=7.0875 PJ=10.8

D039_dim_fail D0_039_dim_fail D1_039_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=8.1 PJ=11.7

D040_dim_fail D0_040_dim_fail D1_040_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.215 PJ=6.3

D041_dim_fail D0_041_dim_fail D1_041_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=2.43 PJ=7.2

D042_dim_fail D0_042_dim_fail D1_042_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=3.645 PJ=8.1

D043_dim_fail D0_043_dim_fail D1_043_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=4.86 PJ=9.0

D044_dim_fail D0_044_dim_fail D1_044_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=6.075 PJ=9.9

D045_dim_fail D0_045_dim_fail D1_045_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=7.29 PJ=10.8

D046_dim_fail D0_046_dim_fail D1_046_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=8.505 PJ=11.7

D047_dim_fail D0_047_dim_fail D1_047_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=9.72 PJ=12.6

D048_dim_fail D0_048_dim_fail D1_048_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.4175 PJ=7.2

D049_dim_fail D0_049_dim_fail D1_049_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=2.835 PJ=8.1

D050_dim_fail D0_050_dim_fail D1_050_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=4.2525 PJ=9.0

D051_dim_fail D0_051_dim_fail D1_051_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=5.67 PJ=9.9

D052_dim_fail D0_052_dim_fail D1_052_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=7.0875 PJ=10.8

D053_dim_fail D0_053_dim_fail D1_053_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=8.505 PJ=11.7

D054_dim_fail D0_054_dim_fail D1_054_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=9.9225 PJ=12.6

D055_dim_fail D0_055_dim_fail D1_055_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=11.34 PJ=13.5

D056_dim_fail D0_056_dim_fail D1_056_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=1.62 PJ=8.1

D057_dim_fail D0_057_dim_fail D1_057_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=3.24 PJ=9.0

D058_dim_fail D0_058_dim_fail D1_058_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=4.86 PJ=9.9

D059_dim_fail D0_059_dim_fail D1_059_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=6.48 PJ=10.8

D060_dim_fail D0_060_dim_fail D1_060_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=8.1 PJ=11.7

D061_dim_fail D0_061_dim_fail D1_061_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=9.72 PJ=12.6

D062_dim_fail D0_062_dim_fail D1_062_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=11.34 PJ=13.5

D063_dim_fail D0_063_dim_fail D1_063_dim_fail sky130_fd_pr__diode_pd2nw_05v5 AREA=12.96 PJ=14.4

.ENDS