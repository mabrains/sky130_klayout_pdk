 
* Copyright 2022 Mabrains
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Affero General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Affero General Public License for more details.
* 
* You should have received a copy of the GNU Affero General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.

.SUBCKT TOP 
+ L0_1 L1_1 TAP_1
+ L0_2 L1_2 TAP_2

X1 L0_1 L1_1 TAP_1 sky130_fd_pr__rf_test_coil1

X2 L0_2 L1_2 TAP_2 sky130_fd_pr__rf_test_coil2

.ENDS

.SUBCKT sky130_fd_pr__rf_test_coil1 L0_1 L1_1 TAP_1

Lx L0_1 L1_1 TAP_1 sky130_fd_pr__rf_ind_03_90

.ENDS

.SUBCKT sky130_fd_pr__rf_test_coil2 L0_2 L1_2 TAP_2

Lx L0_2 L1_2 TAP_2 sky130_fd_pr__rf_ind_05_125

.ENDS


