* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_ls__nand3b_1 A_N B C VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.12U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.12U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.12U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.84U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.74U l=0.15U mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.74U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.74U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.55U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_ls__nand3b_1
