* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_lp__nor4_2 A B C D VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.26U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.26U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.26U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.26U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.84U l=0.15U mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.84U l=0.15U mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.84U l=0.15U mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.84U l=0.15U mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS sky130_fd_sc_lp__nor4_2
