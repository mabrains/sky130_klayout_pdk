* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
*.PININFO DIODE:I VGND:I VNB:I VPB:I VPWR:I
* Notes: Tap diode is not represented here.
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 m=1 A=0.4347p P=2.64u
.ENDS sky130_fd_sc_hd__diode_2
