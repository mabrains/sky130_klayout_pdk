 
* Copyright 2022 Mabrains
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Affero General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Affero General Public License for more details.
* 
* You should have received a copy of the GNU Affero General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM02W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE

Mx_net_fail DRAIN_net_fail GATE_net_fail SOURCE_net_fail SUBSTRATE sky130_fd_pr__rf_nfet_01v8_lvt_bM02W1p65L0p18 w=4.073849999999999u l=0.22221u nf=2 m=1 ad=0.29529239999999995p as=0.29529239999999995p pd=2.752935u ps=2.752935u nrd=0.2170251 nrs=0.2170251 sa=0.0 sb=0.0 sd=0.0

.ENDS