 
* Copyright 2022 Mabrains
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Affero General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Affero General Public License for more details.
* 
* You should have received a copy of the GNU Affero General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.

.SUBCKT sky130_fd_pr__diode_pw2nd_05v5_nvt SUB
+ SUB D1_000
+ SUB D1_001
+ SUB D1_002
+ SUB D1_003
+ SUB D1_004
+ SUB D1_005
+ SUB D1_006
+ SUB D1_007
+ SUB D1_008
+ SUB D1_009
+ SUB D1_010
+ SUB D1_011
+ SUB D1_012
+ SUB D1_013
+ SUB D1_014
+ SUB D1_015
+ SUB D1_016
+ SUB D1_017
+ SUB D1_018
+ SUB D1_019
+ SUB D1_020
+ SUB D1_021
+ SUB D1_022
+ SUB D1_023
+ SUB D1_024
+ SUB D1_025
+ SUB D1_026
+ SUB D1_027
+ SUB D1_028
+ SUB D1_029
+ SUB D1_030
+ SUB D1_031
+ SUB D1_032
+ SUB D1_033
+ SUB D1_034
+ SUB D1_035
+ SUB D1_036
+ SUB D1_037
+ SUB D1_038
+ SUB D1_039
+ SUB D1_040
+ SUB D1_041
+ SUB D1_042
+ SUB D1_043
+ SUB D1_044
+ SUB D1_045
+ SUB D1_046
+ SUB D1_047
+ SUB D1_048
+ SUB D1_049
+ SUB D1_050
+ SUB D1_051
+ SUB D1_052
+ SUB D1_053
+ SUB D1_054
+ SUB D1_055
+ SUB D1_056
+ SUB D1_057
+ SUB D1_058
+ SUB D1_059
+ SUB D1_060
+ SUB D1_061
+ SUB D1_062
+ SUB D1_063

D000 SUB D1_000 sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.2025p P=1.8u

D001 SUB D1_001 sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.405p P=2.7u

D002 SUB D1_002 sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.6075p P=3.6u

D003 SUB D1_003 sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.81p P=4.5u

D004 SUB D1_004 sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.0125p P=5.4u

D005 SUB D1_005 sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.215p P=6.3u

D006 SUB D1_006 sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.4175p P=7.2u

D007 SUB D1_007 sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.62p P=8.1u

D008 SUB D1_008 sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.405p P=2.7u

D009 SUB D1_009 sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.81p P=3.6u

D010 SUB D1_010 sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.215p P=4.5u

D011 SUB D1_011 sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.62p P=5.4u

D012 SUB D1_012 sky130_fd_pr__diode_pw2nd_05v5_nvt A=2.025p P=6.3u

D013 SUB D1_013 sky130_fd_pr__diode_pw2nd_05v5_nvt A=2.43p P=7.2u

D014 SUB D1_014 sky130_fd_pr__diode_pw2nd_05v5_nvt A=2.835p P=8.1u

D015 SUB D1_015 sky130_fd_pr__diode_pw2nd_05v5_nvt A=3.24p P=9.0u

D016 SUB D1_016 sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.6075p P=3.6u

D017 SUB D1_017 sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.215p P=4.5u

D018 SUB D1_018 sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.8225p P=5.4u

D019 SUB D1_019 sky130_fd_pr__diode_pw2nd_05v5_nvt A=2.43p P=6.3u

D020 SUB D1_020 sky130_fd_pr__diode_pw2nd_05v5_nvt A=3.0375p P=7.2u

D021 SUB D1_021 sky130_fd_pr__diode_pw2nd_05v5_nvt A=3.645p P=8.1u

D022 SUB D1_022 sky130_fd_pr__diode_pw2nd_05v5_nvt A=4.2525p P=9.0u

D023 SUB D1_023 sky130_fd_pr__diode_pw2nd_05v5_nvt A=4.86p P=9.9u

D024 SUB D1_024 sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.81p P=4.5u

D025 SUB D1_025 sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.62p P=5.4u

D026 SUB D1_026 sky130_fd_pr__diode_pw2nd_05v5_nvt A=2.43p P=6.3u

D027 SUB D1_027 sky130_fd_pr__diode_pw2nd_05v5_nvt A=3.24p P=7.2u

D028 SUB D1_028 sky130_fd_pr__diode_pw2nd_05v5_nvt A=4.05p P=8.1u

D029 SUB D1_029 sky130_fd_pr__diode_pw2nd_05v5_nvt A=4.86p P=9.0u

D030 SUB D1_030 sky130_fd_pr__diode_pw2nd_05v5_nvt A=5.67p P=9.9u

D031 SUB D1_031 sky130_fd_pr__diode_pw2nd_05v5_nvt A=6.48p P=10.8u

D032 SUB D1_032 sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.0125p P=5.4u

D033 SUB D1_033 sky130_fd_pr__diode_pw2nd_05v5_nvt A=2.025p P=6.3u

D034 SUB D1_034 sky130_fd_pr__diode_pw2nd_05v5_nvt A=3.0375p P=7.2u

D035 SUB D1_035 sky130_fd_pr__diode_pw2nd_05v5_nvt A=4.05p P=8.1u

D036 SUB D1_036 sky130_fd_pr__diode_pw2nd_05v5_nvt A=5.0625p P=9.0u

D037 SUB D1_037 sky130_fd_pr__diode_pw2nd_05v5_nvt A=6.075p P=9.9u

D038 SUB D1_038 sky130_fd_pr__diode_pw2nd_05v5_nvt A=7.0875p P=10.8u

D039 SUB D1_039 sky130_fd_pr__diode_pw2nd_05v5_nvt A=8.1p P=11.7u

D040 SUB D1_040 sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.215p P=6.3u

D041 SUB D1_041 sky130_fd_pr__diode_pw2nd_05v5_nvt A=2.43p P=7.2u

D042 SUB D1_042 sky130_fd_pr__diode_pw2nd_05v5_nvt A=3.645p P=8.1u

D043 SUB D1_043 sky130_fd_pr__diode_pw2nd_05v5_nvt A=4.86p P=9.0u

D044 SUB D1_044 sky130_fd_pr__diode_pw2nd_05v5_nvt A=6.075p P=9.9u

D045 SUB D1_045 sky130_fd_pr__diode_pw2nd_05v5_nvt A=7.29p P=10.8u

D046 SUB D1_046 sky130_fd_pr__diode_pw2nd_05v5_nvt A=8.505p P=11.7u

D047 SUB D1_047 sky130_fd_pr__diode_pw2nd_05v5_nvt A=9.72p P=12.6u

D048 SUB D1_048 sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.4175p P=7.2u

D049 SUB D1_049 sky130_fd_pr__diode_pw2nd_05v5_nvt A=2.835p P=8.1u

D050 SUB D1_050 sky130_fd_pr__diode_pw2nd_05v5_nvt A=4.2525p P=9.0u

D051 SUB D1_051 sky130_fd_pr__diode_pw2nd_05v5_nvt A=5.67p P=9.9u

D052 SUB D1_052 sky130_fd_pr__diode_pw2nd_05v5_nvt A=7.0875p P=10.8u

D053 SUB D1_053 sky130_fd_pr__diode_pw2nd_05v5_nvt A=8.505p P=11.7u

D054 SUB D1_054 sky130_fd_pr__diode_pw2nd_05v5_nvt A=9.9225p P=12.6u

D055 SUB D1_055 sky130_fd_pr__diode_pw2nd_05v5_nvt A=11.34p P=13.5u

D056 SUB D1_056 sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.62p P=8.1u

D057 SUB D1_057 sky130_fd_pr__diode_pw2nd_05v5_nvt A=3.24p P=9.0u

D058 SUB D1_058 sky130_fd_pr__diode_pw2nd_05v5_nvt A=4.86p P=9.9u

D059 SUB D1_059 sky130_fd_pr__diode_pw2nd_05v5_nvt A=6.48p P=10.8u

D060 SUB D1_060 sky130_fd_pr__diode_pw2nd_05v5_nvt A=8.1p P=11.7u

D061 SUB D1_061 sky130_fd_pr__diode_pw2nd_05v5_nvt A=9.72p P=12.6u

D062 SUB D1_062 sky130_fd_pr__diode_pw2nd_05v5_nvt A=11.34p P=13.5u

D063 SUB D1_063 sky130_fd_pr__diode_pw2nd_05v5_nvt A=12.96p P=14.4u

.ENDS