 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8 SUBSTRATE SOURCE0 GATE0 DRAIN0 SOURCE1 GATE1 DRAIN1 SOURCE2 GATE2 DRAIN2 SOURCE3 GATE3 DRAIN3 SOURCE4 GATE4 DRAIN4 SOURCE5 GATE5 DRAIN5 SOURCE6 GATE6 DRAIN6 SOURCE7 GATE7 DRAIN7 SOURCE8 GATE8 DRAIN8 SOURCE9 GATE9 DRAIN9 SOURCE10 GATE10 DRAIN10 SOURCE11 GATE11 DRAIN11 SOURCE12 GATE12 DRAIN12 SOURCE13 GATE13 DRAIN13 SOURCE14 GATE14 DRAIN14 SOURCE15 GATE15 DRAIN15 SOURCE16 GATE16 DRAIN16 SOURCE17 GATE17 DRAIN17 SOURCE18 GATE18 DRAIN18 SOURCE19 GATE19 DRAIN19 SOURCE20 GATE20 DRAIN20 SOURCE21 GATE21 DRAIN21 SOURCE22 GATE22 DRAIN22 SOURCE23 GATE23 DRAIN23 SOURCE24 GATE24 DRAIN24 SOURCE25 GATE25 DRAIN25 SOURCE26 GATE26 DRAIN26 SOURCE27 GATE27 DRAIN27 SOURCE28 GATE28 DRAIN28 SOURCE29 GATE29 DRAIN29 SOURCE30 GATE30 DRAIN30 SOURCE31 GATE31 DRAIN31 SOURCE32 GATE32 DRAIN32 SOURCE33 GATE33 DRAIN33 SOURCE34 GATE34 DRAIN34 SOURCE35 GATE35 DRAIN35 SOURCE36 GATE36 DRAIN36 SOURCE37 GATE37 DRAIN37 SOURCE38 GATE38 DRAIN38 SOURCE39 GATE39 DRAIN39 SOURCE40 GATE40 DRAIN40 SOURCE41 GATE41 DRAIN41 SOURCE42 GATE42 DRAIN42 SOURCE43 GATE43 DRAIN43 SOURCE44 GATE44 DRAIN44 SOURCE45 GATE45 DRAIN45 SOURCE46 GATE46 DRAIN46 SOURCE47 GATE47 DRAIN47 SOURCE48 GATE48 DRAIN48 SOURCE49 GATE49 DRAIN49 SOURCE50 GATE50 DRAIN50 SOURCE51 GATE51 DRAIN51 SOURCE52 GATE52 DRAIN52 SOURCE53 GATE53 DRAIN53 SOURCE54 GATE54 DRAIN54 SOURCE55 GATE55 DRAIN55 SOURCE56 GATE56 DRAIN56 SOURCE57 GATE57 DRAIN57 SOURCE58 GATE58 DRAIN58 SOURCE59 GATE59 DRAIN59 SOURCE60 GATE60 DRAIN60 SOURCE61 GATE61 DRAIN61 SOURCE62 GATE62 DRAIN62 SOURCE63 GATE63 DRAIN63
M0 SOURCE0 GATE0 DRAIN0 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=0.15 nf=1

M1 SOURCE1 GATE1 DRAIN1 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=0.15 nf=1

M2 SOURCE2 GATE2 DRAIN2 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=0.15 nf=1

M3 SOURCE3 GATE3 DRAIN3 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=0.15 nf=1

M4 SOURCE4 GATE4 DRAIN4 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=2.15 nf=1

M5 SOURCE5 GATE5 DRAIN5 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=2.15 nf=1

M6 SOURCE6 GATE6 DRAIN6 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=2.15 nf=1

M7 SOURCE7 GATE7 DRAIN7 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=2.15 nf=1

M8 SOURCE8 GATE8 DRAIN8 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=4.15 nf=1

M9 SOURCE9 GATE9 DRAIN9 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=4.15 nf=1

M10 SOURCE10 GATE10 DRAIN10 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=4.15 nf=1

M11 SOURCE11 GATE11 DRAIN11 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=4.15 nf=1

M12 SOURCE12 GATE12 DRAIN12 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=6.15 nf=1

M13 SOURCE13 GATE13 DRAIN13 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=6.15 nf=1

M14 SOURCE14 GATE14 DRAIN14 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=6.15 nf=1

M15 SOURCE15 GATE15 DRAIN15 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=6.15 nf=1

M16 SOURCE16 GATE16 DRAIN16 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=0.15 nf=5

M17 SOURCE17 GATE17 DRAIN17 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=0.15 nf=5

M18 SOURCE18 GATE18 DRAIN18 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=0.15 nf=5

M19 SOURCE19 GATE19 DRAIN19 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=0.15 nf=5

M20 SOURCE20 GATE20 DRAIN20 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=2.15 nf=5

M21 SOURCE21 GATE21 DRAIN21 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=2.15 nf=5

M22 SOURCE22 GATE22 DRAIN22 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=2.15 nf=5

M23 SOURCE23 GATE23 DRAIN23 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=2.15 nf=5

M24 SOURCE24 GATE24 DRAIN24 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=4.15 nf=5

M25 SOURCE25 GATE25 DRAIN25 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=4.15 nf=5

M26 SOURCE26 GATE26 DRAIN26 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=4.15 nf=5

M27 SOURCE27 GATE27 DRAIN27 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=4.15 nf=5

M28 SOURCE28 GATE28 DRAIN28 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=6.15 nf=5

M29 SOURCE29 GATE29 DRAIN29 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=6.15 nf=5

M30 SOURCE30 GATE30 DRAIN30 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=6.15 nf=5

M31 SOURCE31 GATE31 DRAIN31 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=6.15 nf=5

M32 SOURCE32 GATE32 DRAIN32 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=0.15 nf=9

M33 SOURCE33 GATE33 DRAIN33 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=0.15 nf=9

M34 SOURCE34 GATE34 DRAIN34 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=0.15 nf=9

M35 SOURCE35 GATE35 DRAIN35 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=0.15 nf=9

M36 SOURCE36 GATE36 DRAIN36 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=2.15 nf=9

M37 SOURCE37 GATE37 DRAIN37 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=2.15 nf=9

M38 SOURCE38 GATE38 DRAIN38 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=2.15 nf=9

M39 SOURCE39 GATE39 DRAIN39 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=2.15 nf=9

M40 SOURCE40 GATE40 DRAIN40 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=4.15 nf=9

M41 SOURCE41 GATE41 DRAIN41 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=4.15 nf=9

M42 SOURCE42 GATE42 DRAIN42 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=4.15 nf=9

M43 SOURCE43 GATE43 DRAIN43 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=4.15 nf=9

M44 SOURCE44 GATE44 DRAIN44 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=6.15 nf=9

M45 SOURCE45 GATE45 DRAIN45 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=6.15 nf=9

M46 SOURCE46 GATE46 DRAIN46 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=6.15 nf=9

M47 SOURCE47 GATE47 DRAIN47 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=6.15 nf=9

M48 SOURCE48 GATE48 DRAIN48 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=0.15 nf=13

M49 SOURCE49 GATE49 DRAIN49 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=0.15 nf=13

M50 SOURCE50 GATE50 DRAIN50 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=0.15 nf=13

M51 SOURCE51 GATE51 DRAIN51 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=0.15 nf=13

M52 SOURCE52 GATE52 DRAIN52 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=2.15 nf=13

M53 SOURCE53 GATE53 DRAIN53 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=2.15 nf=13

M54 SOURCE54 GATE54 DRAIN54 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=2.15 nf=13

M55 SOURCE55 GATE55 DRAIN55 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=2.15 nf=13

M56 SOURCE56 GATE56 DRAIN56 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=4.15 nf=13

M57 SOURCE57 GATE57 DRAIN57 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=4.15 nf=13

M58 SOURCE58 GATE58 DRAIN58 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=4.15 nf=13

M59 SOURCE59 GATE59 DRAIN59 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=4.15 nf=13

M60 SOURCE60 GATE60 DRAIN60 SUBSTRATE sky130_fd_pr__nfet_01v8 w=0.42 l=6.15 nf=13

M61 SOURCE61 GATE61 DRAIN61 SUBSTRATE sky130_fd_pr__nfet_01v8 w=2.1 l=6.15 nf=13

M62 SOURCE62 GATE62 DRAIN62 SUBSTRATE sky130_fd_pr__nfet_01v8 w=3.7800000000000002 l=6.15 nf=13

M63 SOURCE63 GATE63 DRAIN63 SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.460000000000001 l=6.15 nf=13

.ENDS