* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_ms__ha_4 A B VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
MMIN2 COUT majb VGND VNB sky130_fd_pr__nfet_01v8_lvt m=4 w=0.74U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB sky130_fd_pr__nfet_01v8_lvt m=4 w=0.74U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB sky130_fd_pr__nfet_01v8_lvt m=2 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB sky130_fd_pr__nfet_01v8_lvt m=2 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB sky130_fd_pr__nfet_01v8_lvt m=2 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB sky130_fd_pr__nfet_01v8_lvt m=2 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB sky130_fd_pr__nfet_01v8_lvt m=2 w=0.64U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB sky130_fd_pr__pfet_01v8 m=4 w=1.12U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB sky130_fd_pr__pfet_01v8 m=4 w=1.12U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB sky130_fd_pr__pfet_01v8 m=2 w=0.84U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB sky130_fd_pr__pfet_01v8 m=2 w=0.84U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB sky130_fd_pr__pfet_01v8 m=2 w=0.84U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8 m=2 w=1.0U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB sky130_fd_pr__pfet_01v8 m=2 w=1.0U l=0.18U mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_ms__ha_4
