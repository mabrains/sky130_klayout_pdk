* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_ls__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMNnor0 inor A1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74U l=0.15U mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12U l=0.15U mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
.ENDS sky130_fd_sc_ls__a2bb2oi_1
