 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__model__cap_mim_m4
+ C0_000 C1_000 C0_000_net_fail C0_000_dim_fail C1_000_net_fail C1_000_dim_fail
+ C0_001 C1_001 C0_001_net_fail C0_001_dim_fail C1_001_net_fail C1_001_dim_fail
+ C0_002 C1_002 C0_002_net_fail C0_002_dim_fail C1_002_net_fail C1_002_dim_fail
+ C0_003 C1_003 C0_003_net_fail C0_003_dim_fail C1_003_net_fail C1_003_dim_fail
+ C0_004 C1_004 C0_004_net_fail C0_004_dim_fail C1_004_net_fail C1_004_dim_fail
+ C0_005 C1_005 C0_005_net_fail C0_005_dim_fail C1_005_net_fail C1_005_dim_fail
+ C0_006 C1_006 C0_006_net_fail C0_006_dim_fail C1_006_net_fail C1_006_dim_fail
+ C0_007 C1_007 C0_007_net_fail C0_007_dim_fail C1_007_net_fail C1_007_dim_fail
+ C0_008 C1_008 C0_008_net_fail C0_008_dim_fail C1_008_net_fail C1_008_dim_fail
+ C0_009 C1_009 C0_009_net_fail C0_009_dim_fail C1_009_net_fail C1_009_dim_fail
+ C0_010 C1_010 C0_010_net_fail C0_010_dim_fail C1_010_net_fail C1_010_dim_fail
+ C0_011 C1_011 C0_011_net_fail C0_011_dim_fail C1_011_net_fail C1_011_dim_fail
+ C0_012 C1_012 C0_012_net_fail C0_012_dim_fail C1_012_net_fail C1_012_dim_fail
+ C0_013 C1_013 C0_013_net_fail C0_013_dim_fail C1_013_net_fail C1_013_dim_fail
+ C0_014 C1_014 C0_014_net_fail C0_014_dim_fail C1_014_net_fail C1_014_dim_fail
+ C0_015 C1_015 C0_015_net_fail C0_015_dim_fail C1_015_net_fail C1_015_dim_fail
+ C0_016 C1_016 C0_016_net_fail C0_016_dim_fail C1_016_net_fail C1_016_dim_fail
+ C0_017 C1_017 C0_017_net_fail C0_017_dim_fail C1_017_net_fail C1_017_dim_fail
+ C0_018 C1_018 C0_018_net_fail C0_018_dim_fail C1_018_net_fail C1_018_dim_fail
+ C0_019 C1_019 C0_019_net_fail C0_019_dim_fail C1_019_net_fail C1_019_dim_fail
+ C0_020 C1_020 C0_020_net_fail C0_020_dim_fail C1_020_net_fail C1_020_dim_fail
+ C0_021 C1_021 C0_021_net_fail C0_021_dim_fail C1_021_net_fail C1_021_dim_fail
+ C0_022 C1_022 C0_022_net_fail C0_022_dim_fail C1_022_net_fail C1_022_dim_fail
+ C0_023 C1_023 C0_023_net_fail C0_023_dim_fail C1_023_net_fail C1_023_dim_fail
+ C0_024 C1_024 C0_024_net_fail C0_024_dim_fail C1_024_net_fail C1_024_dim_fail
+ C0_025 C1_025 C0_025_net_fail C0_025_dim_fail C1_025_net_fail C1_025_dim_fail
+ C0_026 C1_026 C0_026_net_fail C0_026_dim_fail C1_026_net_fail C1_026_dim_fail
+ C0_027 C1_027 C0_027_net_fail C0_027_dim_fail C1_027_net_fail C1_027_dim_fail
+ C0_028 C1_028 C0_028_net_fail C0_028_dim_fail C1_028_net_fail C1_028_dim_fail
+ C0_029 C1_029 C0_029_net_fail C0_029_dim_fail C1_029_net_fail C1_029_dim_fail
+ C0_030 C1_030 C0_030_net_fail C0_030_dim_fail C1_030_net_fail C1_030_dim_fail
+ C0_031 C1_031 C0_031_net_fail C0_031_dim_fail C1_031_net_fail C1_031_dim_fail
+ C0_032 C1_032 C0_032_net_fail C0_032_dim_fail C1_032_net_fail C1_032_dim_fail
+ C0_033 C1_033 C0_033_net_fail C0_033_dim_fail C1_033_net_fail C1_033_dim_fail
+ C0_034 C1_034 C0_034_net_fail C0_034_dim_fail C1_034_net_fail C1_034_dim_fail
+ C0_035 C1_035 C0_035_net_fail C0_035_dim_fail C1_035_net_fail C1_035_dim_fail
+ C0_036 C1_036 C0_036_net_fail C0_036_dim_fail C1_036_net_fail C1_036_dim_fail
+ C0_037 C1_037 C0_037_net_fail C0_037_dim_fail C1_037_net_fail C1_037_dim_fail
+ C0_038 C1_038 C0_038_net_fail C0_038_dim_fail C1_038_net_fail C1_038_dim_fail
+ C0_039 C1_039 C0_039_net_fail C0_039_dim_fail C1_039_net_fail C1_039_dim_fail
+ C0_040 C1_040 C0_040_net_fail C0_040_dim_fail C1_040_net_fail C1_040_dim_fail
+ C0_041 C1_041 C0_041_net_fail C0_041_dim_fail C1_041_net_fail C1_041_dim_fail
+ C0_042 C1_042 C0_042_net_fail C0_042_dim_fail C1_042_net_fail C1_042_dim_fail
+ C0_043 C1_043 C0_043_net_fail C0_043_dim_fail C1_043_net_fail C1_043_dim_fail
+ C0_044 C1_044 C0_044_net_fail C0_044_dim_fail C1_044_net_fail C1_044_dim_fail
+ C0_045 C1_045 C0_045_net_fail C0_045_dim_fail C1_045_net_fail C1_045_dim_fail
+ C0_046 C1_046 C0_046_net_fail C0_046_dim_fail C1_046_net_fail C1_046_dim_fail
+ C0_047 C1_047 C0_047_net_fail C0_047_dim_fail C1_047_net_fail C1_047_dim_fail
+ C0_048 C1_048 C0_048_net_fail C0_048_dim_fail C1_048_net_fail C1_048_dim_fail
+ C0_049 C1_049 C0_049_net_fail C0_049_dim_fail C1_049_net_fail C1_049_dim_fail
+ C0_050 C1_050 C0_050_net_fail C0_050_dim_fail C1_050_net_fail C1_050_dim_fail
+ C0_051 C1_051 C0_051_net_fail C0_051_dim_fail C1_051_net_fail C1_051_dim_fail
+ C0_052 C1_052 C0_052_net_fail C0_052_dim_fail C1_052_net_fail C1_052_dim_fail
+ C0_053 C1_053 C0_053_net_fail C0_053_dim_fail C1_053_net_fail C1_053_dim_fail
+ C0_054 C1_054 C0_054_net_fail C0_054_dim_fail C1_054_net_fail C1_054_dim_fail
+ C0_055 C1_055 C0_055_net_fail C0_055_dim_fail C1_055_net_fail C1_055_dim_fail
+ C0_056 C1_056 C0_056_net_fail C0_056_dim_fail C1_056_net_fail C1_056_dim_fail
+ C0_057 C1_057 C0_057_net_fail C0_057_dim_fail C1_057_net_fail C1_057_dim_fail
+ C0_058 C1_058 C0_058_net_fail C0_058_dim_fail C1_058_net_fail C1_058_dim_fail
+ C0_059 C1_059 C0_059_net_fail C0_059_dim_fail C1_059_net_fail C1_059_dim_fail
+ C0_060 C1_060 C0_060_net_fail C0_060_dim_fail C1_060_net_fail C1_060_dim_fail
+ C0_061 C1_061 C0_061_net_fail C0_061_dim_fail C1_061_net_fail C1_061_dim_fail
+ C0_062 C1_062 C0_062_net_fail C0_062_dim_fail C1_062_net_fail C1_062_dim_fail
+ C0_063 C1_063 C0_063_net_fail C0_063_dim_fail C1_063_net_fail C1_063_dim_fail
+ C0_064 C1_064 C0_064_net_fail C0_064_dim_fail C1_064_net_fail C1_064_dim_fail
+ C0_065 C1_065 C0_065_net_fail C0_065_dim_fail C1_065_net_fail C1_065_dim_fail
+ C0_066 C1_066 C0_066_net_fail C0_066_dim_fail C1_066_net_fail C1_066_dim_fail
+ C0_067 C1_067 C0_067_net_fail C0_067_dim_fail C1_067_net_fail C1_067_dim_fail
+ C0_068 C1_068 C0_068_net_fail C0_068_dim_fail C1_068_net_fail C1_068_dim_fail
+ C0_069 C1_069 C0_069_net_fail C0_069_dim_fail C1_069_net_fail C1_069_dim_fail
+ C0_070 C1_070 C0_070_net_fail C0_070_dim_fail C1_070_net_fail C1_070_dim_fail
+ C0_071 C1_071 C0_071_net_fail C0_071_dim_fail C1_071_net_fail C1_071_dim_fail
+ C0_072 C1_072 C0_072_net_fail C0_072_dim_fail C1_072_net_fail C1_072_dim_fail
+ C0_073 C1_073 C0_073_net_fail C0_073_dim_fail C1_073_net_fail C1_073_dim_fail
+ C0_074 C1_074 C0_074_net_fail C0_074_dim_fail C1_074_net_fail C1_074_dim_fail
+ C0_075 C1_075 C0_075_net_fail C0_075_dim_fail C1_075_net_fail C1_075_dim_fail
+ C0_076 C1_076 C0_076_net_fail C0_076_dim_fail C1_076_net_fail C1_076_dim_fail
+ C0_077 C1_077 C0_077_net_fail C0_077_dim_fail C1_077_net_fail C1_077_dim_fail
+ C0_078 C1_078 C0_078_net_fail C0_078_dim_fail C1_078_net_fail C1_078_dim_fail
+ C0_079 C1_079 C0_079_net_fail C0_079_dim_fail C1_079_net_fail C1_079_dim_fail
+ C0_080 C1_080 C0_080_net_fail C0_080_dim_fail C1_080_net_fail C1_080_dim_fail

C000 C0_000 C1_000 sky130_fd_pr__model__cap_mim_m4 AREA=4 PJ=8

C001 C0_001 C1_001 sky130_fd_pr__model__cap_mim_m4 AREA=24 PJ=28

C002 C0_002 C1_002 sky130_fd_pr__model__cap_mim_m4 AREA=44 PJ=48

C003 C0_003 C1_003 sky130_fd_pr__model__cap_mim_m4 AREA=64 PJ=68

C004 C0_004 C1_004 sky130_fd_pr__model__cap_mim_m4 AREA=84 PJ=88

C005 C0_005 C1_005 sky130_fd_pr__model__cap_mim_m4 AREA=104 PJ=108

C006 C0_006 C1_006 sky130_fd_pr__model__cap_mim_m4 AREA=124 PJ=128

C007 C0_007 C1_007 sky130_fd_pr__model__cap_mim_m4 AREA=144 PJ=148

C008 C0_008 C1_008 sky130_fd_pr__model__cap_mim_m4 AREA=164 PJ=168

C009 C0_009 C1_009 sky130_fd_pr__model__cap_mim_m4 AREA=24 PJ=28

C010 C0_010 C1_010 sky130_fd_pr__model__cap_mim_m4 AREA=144 PJ=48

C011 C0_011 C1_011 sky130_fd_pr__model__cap_mim_m4 AREA=264 PJ=68

C012 C0_012 C1_012 sky130_fd_pr__model__cap_mim_m4 AREA=384 PJ=88

C013 C0_013 C1_013 sky130_fd_pr__model__cap_mim_m4 AREA=504 PJ=108

C014 C0_014 C1_014 sky130_fd_pr__model__cap_mim_m4 AREA=624 PJ=128

C015 C0_015 C1_015 sky130_fd_pr__model__cap_mim_m4 AREA=744 PJ=148

C016 C0_016 C1_016 sky130_fd_pr__model__cap_mim_m4 AREA=864 PJ=168

C017 C0_017 C1_017 sky130_fd_pr__model__cap_mim_m4 AREA=984 PJ=188

C018 C0_018 C1_018 sky130_fd_pr__model__cap_mim_m4 AREA=44 PJ=48

C019 C0_019 C1_019 sky130_fd_pr__model__cap_mim_m4 AREA=264 PJ=68

C020 C0_020 C1_020 sky130_fd_pr__model__cap_mim_m4 AREA=484 PJ=88

C021 C0_021 C1_021 sky130_fd_pr__model__cap_mim_m4 AREA=704 PJ=108

C022 C0_022 C1_022 sky130_fd_pr__model__cap_mim_m4 AREA=924 PJ=128

C023 C0_023 C1_023 sky130_fd_pr__model__cap_mim_m4 AREA=1144 PJ=148

C024 C0_024 C1_024 sky130_fd_pr__model__cap_mim_m4 AREA=1364 PJ=168

C025 C0_025 C1_025 sky130_fd_pr__model__cap_mim_m4 AREA=1584 PJ=188

C026 C0_026 C1_026 sky130_fd_pr__model__cap_mim_m4 AREA=1804 PJ=208

C027 C0_027 C1_027 sky130_fd_pr__model__cap_mim_m4 AREA=64 PJ=68

C028 C0_028 C1_028 sky130_fd_pr__model__cap_mim_m4 AREA=384 PJ=88

C029 C0_029 C1_029 sky130_fd_pr__model__cap_mim_m4 AREA=704 PJ=108

C030 C0_030 C1_030 sky130_fd_pr__model__cap_mim_m4 AREA=1024 PJ=128

C031 C0_031 C1_031 sky130_fd_pr__model__cap_mim_m4 AREA=1344 PJ=148

C032 C0_032 C1_032 sky130_fd_pr__model__cap_mim_m4 AREA=1664 PJ=168

C033 C0_033 C1_033 sky130_fd_pr__model__cap_mim_m4 AREA=1984 PJ=188

C034 C0_034 C1_034 sky130_fd_pr__model__cap_mim_m4 AREA=2304 PJ=208

C035 C0_035 C1_035 sky130_fd_pr__model__cap_mim_m4 AREA=2624 PJ=228

C036 C0_036 C1_036 sky130_fd_pr__model__cap_mim_m4 AREA=84 PJ=88

C037 C0_037 C1_037 sky130_fd_pr__model__cap_mim_m4 AREA=504 PJ=108

C038 C0_038 C1_038 sky130_fd_pr__model__cap_mim_m4 AREA=924 PJ=128

C039 C0_039 C1_039 sky130_fd_pr__model__cap_mim_m4 AREA=1344 PJ=148

C040 C0_040 C1_040 sky130_fd_pr__model__cap_mim_m4 AREA=1764 PJ=168

C041 C0_041 C1_041 sky130_fd_pr__model__cap_mim_m4 AREA=2184 PJ=188

C042 C0_042 C1_042 sky130_fd_pr__model__cap_mim_m4 AREA=2604 PJ=208

C043 C0_043 C1_043 sky130_fd_pr__model__cap_mim_m4 AREA=3024 PJ=228

C044 C0_044 C1_044 sky130_fd_pr__model__cap_mim_m4 AREA=3444 PJ=248

C045 C0_045 C1_045 sky130_fd_pr__model__cap_mim_m4 AREA=104 PJ=108

C046 C0_046 C1_046 sky130_fd_pr__model__cap_mim_m4 AREA=624 PJ=128

C047 C0_047 C1_047 sky130_fd_pr__model__cap_mim_m4 AREA=1144 PJ=148

C048 C0_048 C1_048 sky130_fd_pr__model__cap_mim_m4 AREA=1664 PJ=168

C049 C0_049 C1_049 sky130_fd_pr__model__cap_mim_m4 AREA=2184 PJ=188

C050 C0_050 C1_050 sky130_fd_pr__model__cap_mim_m4 AREA=2704 PJ=208

C051 C0_051 C1_051 sky130_fd_pr__model__cap_mim_m4 AREA=3224 PJ=228

C052 C0_052 C1_052 sky130_fd_pr__model__cap_mim_m4 AREA=3744 PJ=248

C053 C0_053 C1_053 sky130_fd_pr__model__cap_mim_m4 AREA=4264 PJ=268

C054 C0_054 C1_054 sky130_fd_pr__model__cap_mim_m4 AREA=124 PJ=128

C055 C0_055 C1_055 sky130_fd_pr__model__cap_mim_m4 AREA=744 PJ=148

C056 C0_056 C1_056 sky130_fd_pr__model__cap_mim_m4 AREA=1364 PJ=168

C057 C0_057 C1_057 sky130_fd_pr__model__cap_mim_m4 AREA=1984 PJ=188

C058 C0_058 C1_058 sky130_fd_pr__model__cap_mim_m4 AREA=2604 PJ=208

C059 C0_059 C1_059 sky130_fd_pr__model__cap_mim_m4 AREA=3224 PJ=228

C060 C0_060 C1_060 sky130_fd_pr__model__cap_mim_m4 AREA=3844 PJ=248

C061 C0_061 C1_061 sky130_fd_pr__model__cap_mim_m4 AREA=4464 PJ=268

C062 C0_062 C1_062 sky130_fd_pr__model__cap_mim_m4 AREA=5084 PJ=288

C063 C0_063 C1_063 sky130_fd_pr__model__cap_mim_m4 AREA=144 PJ=148

C064 C0_064 C1_064 sky130_fd_pr__model__cap_mim_m4 AREA=864 PJ=168

C065 C0_065 C1_065 sky130_fd_pr__model__cap_mim_m4 AREA=1584 PJ=188

C066 C0_066 C1_066 sky130_fd_pr__model__cap_mim_m4 AREA=2304 PJ=208

C067 C0_067 C1_067 sky130_fd_pr__model__cap_mim_m4 AREA=3024 PJ=228

C068 C0_068 C1_068 sky130_fd_pr__model__cap_mim_m4 AREA=3744 PJ=248

C069 C0_069 C1_069 sky130_fd_pr__model__cap_mim_m4 AREA=4464 PJ=268

C070 C0_070 C1_070 sky130_fd_pr__model__cap_mim_m4 AREA=5184 PJ=288

C071 C0_071 C1_071 sky130_fd_pr__model__cap_mim_m4 AREA=5904 PJ=308

C072 C0_072 C1_072 sky130_fd_pr__model__cap_mim_m4 AREA=164 PJ=168

C073 C0_073 C1_073 sky130_fd_pr__model__cap_mim_m4 AREA=984 PJ=188

C074 C0_074 C1_074 sky130_fd_pr__model__cap_mim_m4 AREA=1804 PJ=208

C075 C0_075 C1_075 sky130_fd_pr__model__cap_mim_m4 AREA=2624 PJ=228

C076 C0_076 C1_076 sky130_fd_pr__model__cap_mim_m4 AREA=3444 PJ=248

C077 C0_077 C1_077 sky130_fd_pr__model__cap_mim_m4 AREA=4264 PJ=268

C078 C0_078 C1_078 sky130_fd_pr__model__cap_mim_m4 AREA=5084 PJ=288

C079 C0_079 C1_079 sky130_fd_pr__model__cap_mim_m4 AREA=5904 PJ=308

C080 C0_080 C1_080 sky130_fd_pr__model__cap_mim_m4 AREA=6724 PJ=328

C000_net_fail C0_000_net_fail C1_000_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=6.0 PJ=12.0

C001_net_fail C0_001_net_fail C1_001_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=36.0 PJ=42.0

C002_net_fail C0_002_net_fail C1_002_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=66.0 PJ=72.0

C003_net_fail C0_003_net_fail C1_003_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=96.0 PJ=102.0

C004_net_fail C0_004_net_fail C1_004_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=126.0 PJ=132.0

C005_net_fail C0_005_net_fail C1_005_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=156.0 PJ=162.0

C006_net_fail C0_006_net_fail C1_006_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=186.0 PJ=192.0

C007_net_fail C0_007_net_fail C1_007_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=216.0 PJ=222.0

C008_net_fail C0_008_net_fail C1_008_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=246.0 PJ=252.0

C009_net_fail C0_009_net_fail C1_009_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=36.0 PJ=42.0

C010_net_fail C0_010_net_fail C1_010_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=216.0 PJ=72.0

C011_net_fail C0_011_net_fail C1_011_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=396.0 PJ=102.0

C012_net_fail C0_012_net_fail C1_012_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=576.0 PJ=132.0

C013_net_fail C0_013_net_fail C1_013_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=756.0 PJ=162.0

C014_net_fail C0_014_net_fail C1_014_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=936.0 PJ=192.0

C015_net_fail C0_015_net_fail C1_015_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=1116.0 PJ=222.0

C016_net_fail C0_016_net_fail C1_016_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=1296.0 PJ=252.0

C017_net_fail C0_017_net_fail C1_017_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=1476.0 PJ=282.0

C018_net_fail C0_018_net_fail C1_018_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=66.0 PJ=72.0

C019_net_fail C0_019_net_fail C1_019_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=396.0 PJ=102.0

C020_net_fail C0_020_net_fail C1_020_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=726.0 PJ=132.0

C021_net_fail C0_021_net_fail C1_021_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=1056.0 PJ=162.0

C022_net_fail C0_022_net_fail C1_022_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=1386.0 PJ=192.0

C023_net_fail C0_023_net_fail C1_023_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=1716.0 PJ=222.0

C024_net_fail C0_024_net_fail C1_024_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=2046.0 PJ=252.0

C025_net_fail C0_025_net_fail C1_025_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=2376.0 PJ=282.0

C026_net_fail C0_026_net_fail C1_026_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=2706.0 PJ=312.0

C027_net_fail C0_027_net_fail C1_027_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=96.0 PJ=102.0

C028_net_fail C0_028_net_fail C1_028_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=576.0 PJ=132.0

C029_net_fail C0_029_net_fail C1_029_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=1056.0 PJ=162.0

C030_net_fail C0_030_net_fail C1_030_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=1536.0 PJ=192.0

C031_net_fail C0_031_net_fail C1_031_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=2016.0 PJ=222.0

C032_net_fail C0_032_net_fail C1_032_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=2496.0 PJ=252.0

C033_net_fail C0_033_net_fail C1_033_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=2976.0 PJ=282.0

C034_net_fail C0_034_net_fail C1_034_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=3456.0 PJ=312.0

C035_net_fail C0_035_net_fail C1_035_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=3936.0 PJ=342.0

C036_net_fail C0_036_net_fail C1_036_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=126.0 PJ=132.0

C037_net_fail C0_037_net_fail C1_037_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=756.0 PJ=162.0

C038_net_fail C0_038_net_fail C1_038_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=1386.0 PJ=192.0

C039_net_fail C0_039_net_fail C1_039_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=2016.0 PJ=222.0

C040_net_fail C0_040_net_fail C1_040_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=2646.0 PJ=252.0

C041_net_fail C0_041_net_fail C1_041_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=3276.0 PJ=282.0

C042_net_fail C0_042_net_fail C1_042_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=3906.0 PJ=312.0

C043_net_fail C0_043_net_fail C1_043_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=4536.0 PJ=342.0

C044_net_fail C0_044_net_fail C1_044_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=5166.0 PJ=372.0

C045_net_fail C0_045_net_fail C1_045_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=156.0 PJ=162.0

C046_net_fail C0_046_net_fail C1_046_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=936.0 PJ=192.0

C047_net_fail C0_047_net_fail C1_047_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=1716.0 PJ=222.0

C048_net_fail C0_048_net_fail C1_048_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=2496.0 PJ=252.0

C049_net_fail C0_049_net_fail C1_049_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=3276.0 PJ=282.0

C050_net_fail C0_050_net_fail C1_050_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=4056.0 PJ=312.0

C051_net_fail C0_051_net_fail C1_051_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=4836.0 PJ=342.0

C052_net_fail C0_052_net_fail C1_052_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=5616.0 PJ=372.0

C053_net_fail C0_053_net_fail C1_053_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=6396.0 PJ=402.0

C054_net_fail C0_054_net_fail C1_054_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=186.0 PJ=192.0

C055_net_fail C0_055_net_fail C1_055_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=1116.0 PJ=222.0

C056_net_fail C0_056_net_fail C1_056_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=2046.0 PJ=252.0

C057_net_fail C0_057_net_fail C1_057_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=2976.0 PJ=282.0

C058_net_fail C0_058_net_fail C1_058_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=3906.0 PJ=312.0

C059_net_fail C0_059_net_fail C1_059_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=4836.0 PJ=342.0

C060_net_fail C0_060_net_fail C1_060_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=5766.0 PJ=372.0

C061_net_fail C0_061_net_fail C1_061_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=6696.0 PJ=402.0

C062_net_fail C0_062_net_fail C1_062_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=7626.0 PJ=432.0

C063_net_fail C0_063_net_fail C1_063_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=216.0 PJ=222.0

C064_net_fail C0_064_net_fail C1_064_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=1296.0 PJ=252.0

C065_net_fail C0_065_net_fail C1_065_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=2376.0 PJ=282.0

C066_net_fail C0_066_net_fail C1_066_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=3456.0 PJ=312.0

C067_net_fail C0_067_net_fail C1_067_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=4536.0 PJ=342.0

C068_net_fail C0_068_net_fail C1_068_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=5616.0 PJ=372.0

C069_net_fail C0_069_net_fail C1_069_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=6696.0 PJ=402.0

C070_net_fail C0_070_net_fail C1_070_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=7776.0 PJ=432.0

C071_net_fail C0_071_net_fail C1_071_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=8856.0 PJ=462.0

C072_net_fail C0_072_net_fail C1_072_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=246.0 PJ=252.0

C073_net_fail C0_073_net_fail C1_073_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=1476.0 PJ=282.0

C074_net_fail C0_074_net_fail C1_074_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=2706.0 PJ=312.0

C075_net_fail C0_075_net_fail C1_075_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=3936.0 PJ=342.0

C076_net_fail C0_076_net_fail C1_076_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=5166.0 PJ=372.0

C077_net_fail C0_077_net_fail C1_077_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=6396.0 PJ=402.0

C078_net_fail C0_078_net_fail C1_078_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=7626.0 PJ=432.0

C079_net_fail C0_079_net_fail C1_079_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=8856.0 PJ=462.0

C080_net_fail C0_080_net_fail C1_080_net_fail sky130_fd_pr__model__cap_mim_m4 AREA=10086.0 PJ=492.0

C000_dim_fail C0_000_dim_fail C1_000_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=4 PJ=8

C001_dim_fail C0_001_dim_fail C1_001_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=24 PJ=28

C002_dim_fail C0_002_dim_fail C1_002_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=44 PJ=48

C003_dim_fail C0_003_dim_fail C1_003_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=64 PJ=68

C004_dim_fail C0_004_dim_fail C1_004_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=84 PJ=88

C005_dim_fail C0_005_dim_fail C1_005_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=104 PJ=108

C006_dim_fail C0_006_dim_fail C1_006_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=124 PJ=128

C007_dim_fail C0_007_dim_fail C1_007_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=144 PJ=148

C008_dim_fail C0_008_dim_fail C1_008_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=164 PJ=168

C009_dim_fail C0_009_dim_fail C1_009_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=24 PJ=28

C010_dim_fail C0_010_dim_fail C1_010_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=144 PJ=48

C011_dim_fail C0_011_dim_fail C1_011_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=264 PJ=68

C012_dim_fail C0_012_dim_fail C1_012_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=384 PJ=88

C013_dim_fail C0_013_dim_fail C1_013_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=504 PJ=108

C014_dim_fail C0_014_dim_fail C1_014_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=624 PJ=128

C015_dim_fail C0_015_dim_fail C1_015_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=744 PJ=148

C016_dim_fail C0_016_dim_fail C1_016_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=864 PJ=168

C017_dim_fail C0_017_dim_fail C1_017_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=984 PJ=188

C018_dim_fail C0_018_dim_fail C1_018_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=44 PJ=48

C019_dim_fail C0_019_dim_fail C1_019_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=264 PJ=68

C020_dim_fail C0_020_dim_fail C1_020_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=484 PJ=88

C021_dim_fail C0_021_dim_fail C1_021_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=704 PJ=108

C022_dim_fail C0_022_dim_fail C1_022_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=924 PJ=128

C023_dim_fail C0_023_dim_fail C1_023_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1144 PJ=148

C024_dim_fail C0_024_dim_fail C1_024_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1364 PJ=168

C025_dim_fail C0_025_dim_fail C1_025_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1584 PJ=188

C026_dim_fail C0_026_dim_fail C1_026_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1804 PJ=208

C027_dim_fail C0_027_dim_fail C1_027_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=64 PJ=68

C028_dim_fail C0_028_dim_fail C1_028_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=384 PJ=88

C029_dim_fail C0_029_dim_fail C1_029_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=704 PJ=108

C030_dim_fail C0_030_dim_fail C1_030_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1024 PJ=128

C031_dim_fail C0_031_dim_fail C1_031_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1344 PJ=148

C032_dim_fail C0_032_dim_fail C1_032_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1664 PJ=168

C033_dim_fail C0_033_dim_fail C1_033_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1984 PJ=188

C034_dim_fail C0_034_dim_fail C1_034_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=2304 PJ=208

C035_dim_fail C0_035_dim_fail C1_035_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=2624 PJ=228

C036_dim_fail C0_036_dim_fail C1_036_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=84 PJ=88

C037_dim_fail C0_037_dim_fail C1_037_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=504 PJ=108

C038_dim_fail C0_038_dim_fail C1_038_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=924 PJ=128

C039_dim_fail C0_039_dim_fail C1_039_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1344 PJ=148

C040_dim_fail C0_040_dim_fail C1_040_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1764 PJ=168

C041_dim_fail C0_041_dim_fail C1_041_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=2184 PJ=188

C042_dim_fail C0_042_dim_fail C1_042_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=2604 PJ=208

C043_dim_fail C0_043_dim_fail C1_043_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=3024 PJ=228

C044_dim_fail C0_044_dim_fail C1_044_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=3444 PJ=248

C045_dim_fail C0_045_dim_fail C1_045_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=104 PJ=108

C046_dim_fail C0_046_dim_fail C1_046_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=624 PJ=128

C047_dim_fail C0_047_dim_fail C1_047_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1144 PJ=148

C048_dim_fail C0_048_dim_fail C1_048_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1664 PJ=168

C049_dim_fail C0_049_dim_fail C1_049_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=2184 PJ=188

C050_dim_fail C0_050_dim_fail C1_050_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=2704 PJ=208

C051_dim_fail C0_051_dim_fail C1_051_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=3224 PJ=228

C052_dim_fail C0_052_dim_fail C1_052_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=3744 PJ=248

C053_dim_fail C0_053_dim_fail C1_053_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=4264 PJ=268

C054_dim_fail C0_054_dim_fail C1_054_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=124 PJ=128

C055_dim_fail C0_055_dim_fail C1_055_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=744 PJ=148

C056_dim_fail C0_056_dim_fail C1_056_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1364 PJ=168

C057_dim_fail C0_057_dim_fail C1_057_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1984 PJ=188

C058_dim_fail C0_058_dim_fail C1_058_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=2604 PJ=208

C059_dim_fail C0_059_dim_fail C1_059_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=3224 PJ=228

C060_dim_fail C0_060_dim_fail C1_060_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=3844 PJ=248

C061_dim_fail C0_061_dim_fail C1_061_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=4464 PJ=268

C062_dim_fail C0_062_dim_fail C1_062_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=5084 PJ=288

C063_dim_fail C0_063_dim_fail C1_063_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=144 PJ=148

C064_dim_fail C0_064_dim_fail C1_064_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=864 PJ=168

C065_dim_fail C0_065_dim_fail C1_065_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1584 PJ=188

C066_dim_fail C0_066_dim_fail C1_066_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=2304 PJ=208

C067_dim_fail C0_067_dim_fail C1_067_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=3024 PJ=228

C068_dim_fail C0_068_dim_fail C1_068_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=3744 PJ=248

C069_dim_fail C0_069_dim_fail C1_069_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=4464 PJ=268

C070_dim_fail C0_070_dim_fail C1_070_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=5184 PJ=288

C071_dim_fail C0_071_dim_fail C1_071_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=5904 PJ=308

C072_dim_fail C0_072_dim_fail C1_072_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=164 PJ=168

C073_dim_fail C0_073_dim_fail C1_073_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=984 PJ=188

C074_dim_fail C0_074_dim_fail C1_074_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=1804 PJ=208

C075_dim_fail C0_075_dim_fail C1_075_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=2624 PJ=228

C076_dim_fail C0_076_dim_fail C1_076_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=3444 PJ=248

C077_dim_fail C0_077_dim_fail C1_077_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=4264 PJ=268

C078_dim_fail C0_078_dim_fail C1_078_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=5084 PJ=288

C079_dim_fail C0_079_dim_fail C1_079_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=5904 PJ=308

C080_dim_fail C0_080_dim_fail C1_080_dim_fail sky130_fd_pr__model__cap_mim_m4 AREA=6724 PJ=328

.ENDS