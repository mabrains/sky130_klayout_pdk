* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https:  www.apache.org licenses LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
*.PININFO A_N:I B_N:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42u l=0.15u mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42u l=0.15u mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42u l=0.15u mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMP3 y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42u l=0.15u mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42u l=0.15u mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42u l=0.15u mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0u l=0.15u mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42u l=0.15u mult=1 sa=0.265 sb=0.265
+ sd=0.28 area=0.063 perim=1.14
MMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42u l=0.15u mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42u l=0.15u mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42u l=0.15u mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42u l=0.15u mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMIN1 B B_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42u l=0.15u mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65u l=0.15u mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
.ENDS sky130_fd_sc_hd__and4bb_1
