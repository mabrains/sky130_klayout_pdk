 
* Copyright 2022 Mabrains
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Affero General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Affero General Public License for more details.
* 
* You should have received a copy of the GNU Affero General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.

.SUBCKT sky130_fd_pr__diode_pw2nd_05v5_nvt 
+ D0_000_net_fail D1_000_net_fail
+ D0_001_net_fail D1_001_net_fail
+ D0_002_net_fail D1_002_net_fail
+ D0_003_net_fail D1_003_net_fail
+ D0_004_net_fail D1_004_net_fail
+ D0_005_net_fail D1_005_net_fail
+ D0_006_net_fail D1_006_net_fail
+ D0_007_net_fail D1_007_net_fail
+ D0_008_net_fail D1_008_net_fail
+ D0_009_net_fail D1_009_net_fail
+ D0_010_net_fail D1_010_net_fail
+ D0_011_net_fail D1_011_net_fail
+ D0_012_net_fail D1_012_net_fail
+ D0_013_net_fail D1_013_net_fail
+ D0_014_net_fail D1_014_net_fail
+ D0_015_net_fail D1_015_net_fail
+ D0_016_net_fail D1_016_net_fail
+ D0_017_net_fail D1_017_net_fail
+ D0_018_net_fail D1_018_net_fail
+ D0_019_net_fail D1_019_net_fail
+ D0_020_net_fail D1_020_net_fail
+ D0_021_net_fail D1_021_net_fail
+ D0_022_net_fail D1_022_net_fail
+ D0_023_net_fail D1_023_net_fail
+ D0_024_net_fail D1_024_net_fail
+ D0_025_net_fail D1_025_net_fail
+ D0_026_net_fail D1_026_net_fail
+ D0_027_net_fail D1_027_net_fail
+ D0_028_net_fail D1_028_net_fail
+ D0_029_net_fail D1_029_net_fail
+ D0_030_net_fail D1_030_net_fail
+ D0_031_net_fail D1_031_net_fail
+ D0_032_net_fail D1_032_net_fail
+ D0_033_net_fail D1_033_net_fail
+ D0_034_net_fail D1_034_net_fail
+ D0_035_net_fail D1_035_net_fail
+ D0_036_net_fail D1_036_net_fail
+ D0_037_net_fail D1_037_net_fail
+ D0_038_net_fail D1_038_net_fail
+ D0_039_net_fail D1_039_net_fail
+ D0_040_net_fail D1_040_net_fail
+ D0_041_net_fail D1_041_net_fail
+ D0_042_net_fail D1_042_net_fail
+ D0_043_net_fail D1_043_net_fail
+ D0_044_net_fail D1_044_net_fail
+ D0_045_net_fail D1_045_net_fail
+ D0_046_net_fail D1_046_net_fail
+ D0_047_net_fail D1_047_net_fail
+ D0_048_net_fail D1_048_net_fail
+ D0_049_net_fail D1_049_net_fail
+ D0_050_net_fail D1_050_net_fail
+ D0_051_net_fail D1_051_net_fail
+ D0_052_net_fail D1_052_net_fail
+ D0_053_net_fail D1_053_net_fail
+ D0_054_net_fail D1_054_net_fail
+ D0_055_net_fail D1_055_net_fail
+ D0_056_net_fail D1_056_net_fail
+ D0_057_net_fail D1_057_net_fail
+ D0_058_net_fail D1_058_net_fail
+ D0_059_net_fail D1_059_net_fail
+ D0_060_net_fail D1_060_net_fail
+ D0_061_net_fail D1_061_net_fail
+ D0_062_net_fail D1_062_net_fail
+ D0_063_net_fail D1_063_net_fail

D000_net_fail D0_000_net_fail D1_000_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.24998625p P=2.2220999999999997u

D001_net_fail D0_001_net_fail D1_001_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.4999725p P=3.33315u

D002_net_fail D0_002_net_fail D1_002_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.74995875p P=4.4441999999999995u

D003_net_fail D0_003_net_fail D1_003_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.999945p P=5.55525u

D004_net_fail D0_004_net_fail D1_004_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.24993125p P=6.6663u

D005_net_fail D0_005_net_fail D1_005_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.4999175p P=7.777349999999999u

D006_net_fail D0_006_net_fail D1_006_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.7499037499999999p P=8.888399999999999u

D007_net_fail D0_007_net_fail D1_007_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.99989p P=9.99945u

D008_net_fail D0_008_net_fail D1_008_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.4999725p P=3.33315u

D009_net_fail D0_009_net_fail D1_009_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.999945p P=4.4441999999999995u

D010_net_fail D0_010_net_fail D1_010_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.4999175p P=5.55525u

D011_net_fail D0_011_net_fail D1_011_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.99989p P=6.6663u

D012_net_fail D0_012_net_fail D1_012_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=2.4998625p P=7.777349999999999u

D013_net_fail D0_013_net_fail D1_013_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=2.999835p P=8.888399999999999u

D014_net_fail D0_014_net_fail D1_014_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=3.4998074999999997p P=9.99945u

D015_net_fail D0_015_net_fail D1_015_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=3.99978p P=11.1105u

D016_net_fail D0_016_net_fail D1_016_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.74995875p P=4.4441999999999995u

D017_net_fail D0_017_net_fail D1_017_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.4999175p P=5.55525u

D018_net_fail D0_018_net_fail D1_018_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=2.24987625p P=6.6663u

D019_net_fail D0_019_net_fail D1_019_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=2.999835p P=7.777349999999999u

D020_net_fail D0_020_net_fail D1_020_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=3.74979375p P=8.888399999999999u

D021_net_fail D0_021_net_fail D1_021_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=4.4997525p P=9.99945u

D022_net_fail D0_022_net_fail D1_022_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=5.24971125p P=11.1105u

D023_net_fail D0_023_net_fail D1_023_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=5.99967p P=12.22155u

D024_net_fail D0_024_net_fail D1_024_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=0.999945p P=5.55525u

D025_net_fail D0_025_net_fail D1_025_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.99989p P=6.6663u

D026_net_fail D0_026_net_fail D1_026_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=2.999835p P=7.777349999999999u

D027_net_fail D0_027_net_fail D1_027_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=3.99978p P=8.888399999999999u

D028_net_fail D0_028_net_fail D1_028_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=4.999725p P=9.99945u

D029_net_fail D0_029_net_fail D1_029_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=5.99967p P=11.1105u

D030_net_fail D0_030_net_fail D1_030_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=6.9996149999999995p P=12.22155u

D031_net_fail D0_031_net_fail D1_031_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=7.99956p P=13.3326u

D032_net_fail D0_032_net_fail D1_032_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.24993125p P=6.6663u

D033_net_fail D0_033_net_fail D1_033_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=2.4998625p P=7.777349999999999u

D034_net_fail D0_034_net_fail D1_034_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=3.74979375p P=8.888399999999999u

D035_net_fail D0_035_net_fail D1_035_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=4.999725p P=9.99945u

D036_net_fail D0_036_net_fail D1_036_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=6.249656249999999p P=11.1105u

D037_net_fail D0_037_net_fail D1_037_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=7.4995875p P=12.22155u

D038_net_fail D0_038_net_fail D1_038_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=8.74951875p P=13.3326u

D039_net_fail D0_039_net_fail D1_039_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=9.99945p P=14.443649999999998u

D040_net_fail D0_040_net_fail D1_040_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.4999175p P=7.777349999999999u

D041_net_fail D0_041_net_fail D1_041_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=2.999835p P=8.888399999999999u

D042_net_fail D0_042_net_fail D1_042_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=4.4997525p P=9.99945u

D043_net_fail D0_043_net_fail D1_043_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=5.99967p P=11.1105u

D044_net_fail D0_044_net_fail D1_044_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=7.4995875p P=12.22155u

D045_net_fail D0_045_net_fail D1_045_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=8.999505p P=13.3326u

D046_net_fail D0_046_net_fail D1_046_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=10.4994225p P=14.443649999999998u

D047_net_fail D0_047_net_fail D1_047_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=11.99934p P=15.554699999999999u

D048_net_fail D0_048_net_fail D1_048_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.7499037499999999p P=8.888399999999999u

D049_net_fail D0_049_net_fail D1_049_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=3.4998074999999997p P=9.99945u

D050_net_fail D0_050_net_fail D1_050_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=5.24971125p P=11.1105u

D051_net_fail D0_051_net_fail D1_051_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=6.9996149999999995p P=12.22155u

D052_net_fail D0_052_net_fail D1_052_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=8.74951875p P=13.3326u

D053_net_fail D0_053_net_fail D1_053_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=10.4994225p P=14.443649999999998u

D054_net_fail D0_054_net_fail D1_054_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=12.24932625p P=15.554699999999999u

D055_net_fail D0_055_net_fail D1_055_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=13.999229999999999p P=16.66575u

D056_net_fail D0_056_net_fail D1_056_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=1.99989p P=9.99945u

D057_net_fail D0_057_net_fail D1_057_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=3.99978p P=11.1105u

D058_net_fail D0_058_net_fail D1_058_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=5.99967p P=12.22155u

D059_net_fail D0_059_net_fail D1_059_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=7.99956p P=13.3326u

D060_net_fail D0_060_net_fail D1_060_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=9.99945p P=14.443649999999998u

D061_net_fail D0_061_net_fail D1_061_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=11.99934p P=15.554699999999999u

D062_net_fail D0_062_net_fail D1_062_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=13.999229999999999p P=16.66575u

D063_net_fail D0_063_net_fail D1_063_net_fail sky130_fd_pr__diode_pw2nd_05v5_nvt A=15.99912p P=17.776799999999998u

.ENDS