 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_22p5x23p1_pol1m1m2m3m4m5_noshield 

Cx  sky130_fd_pr__cap_vpp_22p5x23p1_pol1m1m2m3m4m5_noshield

Cx_net_fail  sky130_fd_pr__cap_vpp_22p5x23p1_pol1m1m2m3m4m5_noshield

Cx_dim_fail  sky130_fd_pr__cap_vpp_22p5x23p1_pol1m1m2m3m4m5_noshield

.ENDS