* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4 VPWR A X VPWRIN VPB VGND
M0 a_1032_911 a_620_911 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=0.79u l=0.15u
M1 VPWR a_1032_911 X VPB sky130_fd_pr__pfet_01v8_hvt w=1u l=0.15u M=4
M2 VGND A a_714_47 VGND sky130_fd_pr__nfet_01v8 w=0.65u l=0.15u M=4
M3 VGND a_505_297 a_620_911 VGND sky130_fd_pr__nfet_01v8 w=0.65u l=0.15u M=4
M4 X a_1032_911 VGND VGND sky130_fd_pr__nfet_01v8 w=0.65u l=0.15u M=4
M5 a_1032_911 a_620_911 VGND VGND sky130_fd_pr__nfet_01v8 w=0.65u l=0.15u
M6 a_505_297 A VPWRIN VPWRIN sky130_fd_pr__pfet_01v8_hvt w=1u l=0.15u
M7 VPWR a_714_47 a_620_911 VPB sky130_fd_pr__pfet_01v8_hvt w=0.79u l=0.15u
M8 VPWR a_620_911 a_714_47 VPB sky130_fd_pr__pfet_01v8_hvt w=0.79u l=0.15u
M9 a_505_297 A VGND VGND sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
.ends

