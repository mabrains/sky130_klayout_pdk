* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https:  www.apache.org licenses LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_12 KAPWR VGND VNB VPB VPWR
*.PININFO KAPWR:I VGND:I VNB:I VPB:I VPWR:I
MI1 VGND KAPWR VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55u l=4.73u mult=1 sa=0.265
+ sb=0.265 sd=0.28 area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.87u l=4.73u mult=1
+ sa=0.265 sb=0.265 sd=0.28 area=0.063 perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_decapkapwr_12
