 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT cap_var SUBSTRATE
+ C0_000 C1_000
+ C0_031 C1_031
+ C0_063 C1_063
+ C0_000 C1_000
+ C0_031 C1_031
+ C0_063 C1_063


C000 C0_000 C1_000 SUBSTRATE sky130_fd_pr__cap_var_hvt w=1 l=0.18 nf=1

C031 C0_031 C1_031 SUBSTRATE sky130_fd_pr__cap_var_hvt w=4 l=0.72 nf=5

C063 C0_063 C1_063 SUBSTRATE sky130_fd_pr__cap_var_hvt w=4 l=0.72 nf=13

C000 C0_000 C1_000 SUBSTRATE sky130_fd_pr__cap_var_lvt w=1 l=0.18 nf=1

C031 C0_031 C1_031 SUBSTRATE sky130_fd_pr__cap_var_lvt w=4 l=0.72 nf=5

C063 C0_063 C1_063 SUBSTRATE sky130_fd_pr__cap_var_lvt w=4 l=0.72 nf=13

.ENDS