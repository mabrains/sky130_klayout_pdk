 
* Copyright 2022 Mabrains
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Affero General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Affero General Public License for more details.
* 
* You should have received a copy of the GNU Affero General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.

.SUBCKT sky130_fd_pr__res_xhigh_po_0p69 
+ R0_000_dim_fail R1_000_dim_fail
+ R0_001_dim_fail R1_001_dim_fail
+ R0_002_dim_fail R1_002_dim_fail
+ R0_003_dim_fail R1_003_dim_fail
+ R0_004_dim_fail R1_004_dim_fail
+ R0_005_dim_fail R1_005_dim_fail
+ R0_006_dim_fail R1_006_dim_fail
+ R0_007_dim_fail R1_007_dim_fail
+ R0_008_dim_fail R1_008_dim_fail
+ R0_009_dim_fail R1_009_dim_fail
+ R0_010_dim_fail R1_010_dim_fail
+ R0_011_dim_fail R1_011_dim_fail
+ R0_012_dim_fail R1_012_dim_fail
+ R0_013_dim_fail R1_013_dim_fail
+ R0_014_dim_fail R1_014_dim_fail
+ R0_015_dim_fail R1_015_dim_fail
+ R0_016_dim_fail R1_016_dim_fail
+ R0_017_dim_fail R1_017_dim_fail
+ R0_018_dim_fail R1_018_dim_fail
+ R0_019_dim_fail R1_019_dim_fail
+ R0_020_dim_fail R1_020_dim_fail
+ R0_021_dim_fail R1_021_dim_fail
+ R0_022_dim_fail R1_022_dim_fail
+ R0_023_dim_fail R1_023_dim_fail
+ R0_024_dim_fail R1_024_dim_fail
+ R0_025_dim_fail R1_025_dim_fail
+ R0_026_dim_fail R1_026_dim_fail
+ R0_027_dim_fail R1_027_dim_fail
+ R0_028_dim_fail R1_028_dim_fail
+ R0_029_dim_fail R1_029_dim_fail
+ R0_030_dim_fail R1_030_dim_fail
+ R0_031_dim_fail R1_031_dim_fail
+ R0_032_dim_fail R1_032_dim_fail
+ R0_033_dim_fail R1_033_dim_fail
+ R0_034_dim_fail R1_034_dim_fail
+ R0_035_dim_fail R1_035_dim_fail
+ R0_036_dim_fail R1_036_dim_fail
+ R0_037_dim_fail R1_037_dim_fail
+ R0_038_dim_fail R1_038_dim_fail
+ R0_039_dim_fail R1_039_dim_fail
+ R0_040_dim_fail R1_040_dim_fail
+ R0_041_dim_fail R1_041_dim_fail
+ R0_042_dim_fail R1_042_dim_fail
+ R0_043_dim_fail R1_043_dim_fail
+ R0_044_dim_fail R1_044_dim_fail
+ R0_045_dim_fail R1_045_dim_fail
+ R0_046_dim_fail R1_046_dim_fail
+ R0_047_dim_fail R1_047_dim_fail
+ R0_048_dim_fail R1_048_dim_fail
+ R0_049_dim_fail R1_049_dim_fail
+ R0_050_dim_fail R1_050_dim_fail
+ R0_051_dim_fail R1_051_dim_fail
+ R0_052_dim_fail R1_052_dim_fail
+ R0_053_dim_fail R1_053_dim_fail
+ R0_054_dim_fail R1_054_dim_fail
+ R0_055_dim_fail R1_055_dim_fail
+ R0_056_dim_fail R1_056_dim_fail
+ R0_057_dim_fail R1_057_dim_fail
+ R0_058_dim_fail R1_058_dim_fail
+ R0_059_dim_fail R1_059_dim_fail
+ R0_060_dim_fail R1_060_dim_fail
+ R0_061_dim_fail R1_061_dim_fail
+ R0_062_dim_fail R1_062_dim_fail
+ R0_063_dim_fail R1_063_dim_fail

R000_dim_fail R0_000_dim_fail R1_000_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=1.19u w=0.69u

R001_dim_fail R0_001_dim_fail R1_001_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=2.38u w=0.69u

R002_dim_fail R0_002_dim_fail R1_002_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=3.57u w=0.69u

R003_dim_fail R0_003_dim_fail R1_003_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=4.76u w=0.69u

R004_dim_fail R0_004_dim_fail R1_004_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=5.95u w=0.69u

R005_dim_fail R0_005_dim_fail R1_005_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=7.14u w=0.69u

R006_dim_fail R0_006_dim_fail R1_006_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=8.33u w=0.69u

R007_dim_fail R0_007_dim_fail R1_007_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=9.52u w=0.69u

R008_dim_fail R0_008_dim_fail R1_008_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=2.38u w=0.69u

R009_dim_fail R0_009_dim_fail R1_009_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=4.76u w=0.69u

R010_dim_fail R0_010_dim_fail R1_010_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=7.14u w=0.69u

R011_dim_fail R0_011_dim_fail R1_011_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=9.52u w=0.69u

R012_dim_fail R0_012_dim_fail R1_012_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=11.9u w=0.69u

R013_dim_fail R0_013_dim_fail R1_013_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=14.28u w=0.69u

R014_dim_fail R0_014_dim_fail R1_014_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=16.66u w=0.69u

R015_dim_fail R0_015_dim_fail R1_015_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=19.04u w=0.69u

R016_dim_fail R0_016_dim_fail R1_016_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=3.57u w=0.69u

R017_dim_fail R0_017_dim_fail R1_017_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=7.14u w=0.69u

R018_dim_fail R0_018_dim_fail R1_018_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=10.71u w=0.69u

R019_dim_fail R0_019_dim_fail R1_019_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=14.28u w=0.69u

R020_dim_fail R0_020_dim_fail R1_020_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=17.85u w=0.69u

R021_dim_fail R0_021_dim_fail R1_021_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=21.42u w=0.69u

R022_dim_fail R0_022_dim_fail R1_022_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=24.99u w=0.69u

R023_dim_fail R0_023_dim_fail R1_023_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=28.56u w=0.69u

R024_dim_fail R0_024_dim_fail R1_024_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=4.76u w=0.69u

R025_dim_fail R0_025_dim_fail R1_025_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=9.52u w=0.69u

R026_dim_fail R0_026_dim_fail R1_026_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=14.28u w=0.69u

R027_dim_fail R0_027_dim_fail R1_027_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=19.04u w=0.69u

R028_dim_fail R0_028_dim_fail R1_028_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=23.8u w=0.69u

R029_dim_fail R0_029_dim_fail R1_029_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=28.56u w=0.69u

R030_dim_fail R0_030_dim_fail R1_030_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=33.32u w=0.69u

R031_dim_fail R0_031_dim_fail R1_031_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=38.08u w=0.69u

R032_dim_fail R0_032_dim_fail R1_032_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=5.95u w=0.69u

R033_dim_fail R0_033_dim_fail R1_033_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=11.9u w=0.69u

R034_dim_fail R0_034_dim_fail R1_034_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=17.85u w=0.69u

R035_dim_fail R0_035_dim_fail R1_035_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=23.8u w=0.69u

R036_dim_fail R0_036_dim_fail R1_036_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=29.75u w=0.69u

R037_dim_fail R0_037_dim_fail R1_037_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=35.7u w=0.69u

R038_dim_fail R0_038_dim_fail R1_038_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=41.65u w=0.69u

R039_dim_fail R0_039_dim_fail R1_039_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=47.6u w=0.69u

R040_dim_fail R0_040_dim_fail R1_040_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=7.14u w=0.69u

R041_dim_fail R0_041_dim_fail R1_041_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=14.28u w=0.69u

R042_dim_fail R0_042_dim_fail R1_042_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=21.42u w=0.69u

R043_dim_fail R0_043_dim_fail R1_043_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=28.56u w=0.69u

R044_dim_fail R0_044_dim_fail R1_044_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=35.7u w=0.69u

R045_dim_fail R0_045_dim_fail R1_045_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=42.84u w=0.69u

R046_dim_fail R0_046_dim_fail R1_046_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=49.98u w=0.69u

R047_dim_fail R0_047_dim_fail R1_047_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=57.12u w=0.69u

R048_dim_fail R0_048_dim_fail R1_048_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=8.33u w=0.69u

R049_dim_fail R0_049_dim_fail R1_049_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=16.66u w=0.69u

R050_dim_fail R0_050_dim_fail R1_050_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=24.99u w=0.69u

R051_dim_fail R0_051_dim_fail R1_051_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=33.32u w=0.69u

R052_dim_fail R0_052_dim_fail R1_052_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=41.65u w=0.69u

R053_dim_fail R0_053_dim_fail R1_053_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=49.98u w=0.69u

R054_dim_fail R0_054_dim_fail R1_054_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=58.31u w=0.69u

R055_dim_fail R0_055_dim_fail R1_055_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=66.64u w=0.69u

R056_dim_fail R0_056_dim_fail R1_056_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=9.52u w=0.69u

R057_dim_fail R0_057_dim_fail R1_057_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=19.04u w=0.69u

R058_dim_fail R0_058_dim_fail R1_058_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=28.56u w=0.69u

R059_dim_fail R0_059_dim_fail R1_059_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=38.08u w=0.69u

R060_dim_fail R0_060_dim_fail R1_060_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=47.6u w=0.69u

R061_dim_fail R0_061_dim_fail R1_061_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=57.12u w=0.69u

R062_dim_fail R0_062_dim_fail R1_062_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=66.64u w=0.69u

R063_dim_fail R0_063_dim_fail R1_063_dim_fail sky130_fd_pr__res_xhigh_po_0p69 l=76.16u w=0.69u

.ENDS