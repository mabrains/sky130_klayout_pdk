 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_mcM04W5p00L0p15 Bulk DRAIN GATE SOURCE

Mx Bulk DRAIN GATE SOURCE sky130_fd_pr__rf_pfet_01v8_mcM04W5p00L0p15

Mx_net_fail Bulk_net_fail DRAIN_net_fail GATE_net_fail SOURCE_net_fail sky130_fd_pr__rf_pfet_01v8_mcM04W5p00L0p15

Mx_dim_fail Bulk_dim_fail DRAIN_dim_fail GATE_dim_fail SOURCE_dim_fail sky130_fd_pr__rf_pfet_01v8_mcM04W5p00L0p15

.ENDS