 
# Copyright 2022 SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_aura_blocking B_P D_N2 D_P D_P2 G G_N2 G_P G_P2 NWELL S S_N2 S_P S_P2 VGND VPWR

Xx B_P D_N2 D_P D_P2 G G_N2 G_P G_P2 NWELL S S_N2 S_P S_P2 VGND VPWR sky130_fd_pr__rf_aura_blocking

.ENDS 
